LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.parameters.ALL;

  ENTITY  top IS
  GENERIC (
    BITS : NATURAL := BITS;
    NUM_INPUTS : NATURAL := 784;
    TOTAL_BITS : NATURAL := 6272
  );
  PORT (
      clk, rst, update_weights: IN STD_LOGIC;
      IO_in: IN signed(TOTAL_BITS - 1 DOWNTO 0);
      c0_n0_W_in, c0_n1_W_in, c0_n2_W_in, c0_n3_W_in, c0_n4_W_in, c0_n5_W_in, c0_n6_W_in, c0_n7_W_in, c0_n8_W_in, c0_n9_W_in, c0_n10_W_in, c0_n11_W_in, c0_n12_W_in, c0_n13_W_in, c0_n14_W_in, c0_n15_W_in, c0_n16_W_in, c0_n17_W_in, c0_n18_W_in, c0_n19_W_in, c0_n20_W_in, c0_n21_W_in, c0_n22_W_in, c0_n23_W_in, c0_n24_W_in, c0_n25_W_in, c0_n26_W_in, c0_n27_W_in, c0_n28_W_in, c0_n29_W_in, c0_n30_W_in, c0_n31_W_in, c0_n32_W_in, c0_n33_W_in, c0_n34_W_in, c0_n35_W_in, c0_n36_W_in, c0_n37_W_in, c0_n38_W_in, c0_n39_W_in, c0_n40_W_in, c0_n41_W_in, c0_n42_W_in, c0_n43_W_in, c0_n44_W_in, c0_n45_W_in, c0_n46_W_in, c0_n47_W_in, c0_n48_W_in, c0_n49_W_in, c0_n50_W_in, c0_n51_W_in, c0_n52_W_in, c0_n53_W_in, c0_n54_W_in, c0_n55_W_in, c0_n56_W_in, c0_n57_W_in, c0_n58_W_in, c0_n59_W_in, c0_n60_W_in, c0_n61_W_in, c0_n62_W_in, c0_n63_W_in, c0_n64_W_in, c0_n65_W_in, c0_n66_W_in, c0_n67_W_in, c0_n68_W_in, c0_n69_W_in, c0_n70_W_in, c0_n71_W_in, c0_n72_W_in, c0_n73_W_in, c0_n74_W_in, c0_n75_W_in, c0_n76_W_in, c0_n77_W_in, c0_n78_W_in, c0_n79_W_in, c0_n80_W_in, c0_n81_W_in, c0_n82_W_in, c0_n83_W_in, c0_n84_W_in, c0_n85_W_in, c0_n86_W_in, c0_n87_W_in, c0_n88_W_in, c0_n89_W_in, c0_n90_W_in, c0_n91_W_in, c0_n92_W_in, c0_n93_W_in, c0_n94_W_in, c0_n95_W_in, c0_n96_W_in, c0_n97_W_in, c0_n98_W_in, c0_n99_W_in, c0_n100_W_in, c0_n101_W_in, c0_n102_W_in, c0_n103_W_in, c0_n104_W_in, c0_n105_W_in, c0_n106_W_in, c0_n107_W_in, c0_n108_W_in, c0_n109_W_in, c0_n110_W_in, c0_n111_W_in, c0_n112_W_in, c0_n113_W_in, c0_n114_W_in, c0_n115_W_in, c0_n116_W_in, c0_n117_W_in, c0_n118_W_in, c0_n119_W_in, c0_n120_W_in, c0_n121_W_in, c0_n122_W_in, c0_n123_W_in, c0_n124_W_in, c0_n125_W_in, c0_n126_W_in, c0_n127_W_in, c0_n128_W_in, c0_n129_W_in, c0_n130_W_in, c0_n131_W_in, c0_n132_W_in, c0_n133_W_in, c0_n134_W_in, c0_n135_W_in, c0_n136_W_in, c0_n137_W_in, c0_n138_W_in, c0_n139_W_in, c0_n140_W_in, c0_n141_W_in, c0_n142_W_in, c0_n143_W_in, c0_n144_W_in, c0_n145_W_in, c0_n146_W_in, c0_n147_W_in, c0_n148_W_in, c0_n149_W_in, c0_n150_W_in, c0_n151_W_in, c0_n152_W_in, c0_n153_W_in, c0_n154_W_in, c0_n155_W_in, c0_n156_W_in, c0_n157_W_in, c0_n158_W_in, c0_n159_W_in, c0_n160_W_in, c0_n161_W_in, c0_n162_W_in, c0_n163_W_in, c0_n164_W_in, c0_n165_W_in, c0_n166_W_in, c0_n167_W_in, c0_n168_W_in, c0_n169_W_in, c0_n170_W_in, c0_n171_W_in, c0_n172_W_in, c0_n173_W_in, c0_n174_W_in, c0_n175_W_in, c0_n176_W_in, c0_n177_W_in, c0_n178_W_in, c0_n179_W_in, c0_n180_W_in, c0_n181_W_in, c0_n182_W_in, c0_n183_W_in, c0_n184_W_in, c0_n185_W_in, c0_n186_W_in, c0_n187_W_in, c0_n188_W_in, c0_n189_W_in, c0_n190_W_in, c0_n191_W_in, c0_n192_W_in, c0_n193_W_in, c0_n194_W_in, c0_n195_W_in, c0_n196_W_in, c0_n197_W_in, c0_n198_W_in, c0_n199_W_in, c0_n200_W_in, c0_n201_W_in, c0_n202_W_in, c0_n203_W_in, c0_n204_W_in, c0_n205_W_in, c0_n206_W_in, c0_n207_W_in, c0_n208_W_in, c0_n209_W_in, c0_n210_W_in, c0_n211_W_in, c0_n212_W_in, c0_n213_W_in, c0_n214_W_in, c0_n215_W_in, c0_n216_W_in, c0_n217_W_in, c0_n218_W_in, c0_n219_W_in, c0_n220_W_in, c0_n221_W_in, c0_n222_W_in, c0_n223_W_in, c0_n224_W_in, c0_n225_W_in, c0_n226_W_in, c0_n227_W_in, c0_n228_W_in, c0_n229_W_in, c0_n230_W_in, c0_n231_W_in, c0_n232_W_in, c0_n233_W_in, c0_n234_W_in, c0_n235_W_in, c0_n236_W_in, c0_n237_W_in, c0_n238_W_in, c0_n239_W_in, c0_n240_W_in, c0_n241_W_in, c0_n242_W_in, c0_n243_W_in, c0_n244_W_in, c0_n245_W_in, c0_n246_W_in, c0_n247_W_in, c0_n248_W_in, c0_n249_W_in, c0_n250_W_in, c0_n251_W_in, c0_n252_W_in, c0_n253_W_in, c0_n254_W_in, c0_n255_W_in, c0_n256_W_in, c0_n257_W_in, c0_n258_W_in, c0_n259_W_in, c0_n260_W_in, c0_n261_W_in, c0_n262_W_in, c0_n263_W_in, c0_n264_W_in, c0_n265_W_in, c0_n266_W_in, c0_n267_W_in, c0_n268_W_in, c0_n269_W_in, c0_n270_W_in, c0_n271_W_in, c0_n272_W_in, c0_n273_W_in, c0_n274_W_in, c0_n275_W_in, c0_n276_W_in, c0_n277_W_in, c0_n278_W_in, c0_n279_W_in, c0_n280_W_in, c0_n281_W_in, c0_n282_W_in, c0_n283_W_in, c0_n284_W_in, c0_n285_W_in, c0_n286_W_in, c0_n287_W_in, c0_n288_W_in, c0_n289_W_in, c0_n290_W_in, c0_n291_W_in, c0_n292_W_in, c0_n293_W_in, c0_n294_W_in, c0_n295_W_in, c0_n296_W_in, c0_n297_W_in, c0_n298_W_in, c0_n299_W_in, c0_n300_W_in, c0_n301_W_in, c0_n302_W_in, c0_n303_W_in, c0_n304_W_in, c0_n305_W_in, c0_n306_W_in, c0_n307_W_in, c0_n308_W_in, c0_n309_W_in, c0_n310_W_in, c0_n311_W_in, c0_n312_W_in, c0_n313_W_in, c0_n314_W_in, c0_n315_W_in, c0_n316_W_in, c0_n317_W_in, c0_n318_W_in, c0_n319_W_in, c0_n320_W_in, c0_n321_W_in, c0_n322_W_in, c0_n323_W_in, c0_n324_W_in, c0_n325_W_in, c0_n326_W_in, c0_n327_W_in, c0_n328_W_in, c0_n329_W_in, c0_n330_W_in, c0_n331_W_in, c0_n332_W_in, c0_n333_W_in, c0_n334_W_in, c0_n335_W_in, c0_n336_W_in, c0_n337_W_in, c0_n338_W_in, c0_n339_W_in, c0_n340_W_in, c0_n341_W_in, c0_n342_W_in, c0_n343_W_in, c0_n344_W_in, c0_n345_W_in, c0_n346_W_in, c0_n347_W_in, c0_n348_W_in, c0_n349_W_in, c0_n350_W_in, c0_n351_W_in, c0_n352_W_in, c0_n353_W_in, c0_n354_W_in, c0_n355_W_in, c0_n356_W_in, c0_n357_W_in, c0_n358_W_in, c0_n359_W_in, c0_n360_W_in, c0_n361_W_in, c0_n362_W_in, c0_n363_W_in, c0_n364_W_in, c0_n365_W_in, c0_n366_W_in, c0_n367_W_in, c0_n368_W_in, c0_n369_W_in, c0_n370_W_in, c0_n371_W_in, c0_n372_W_in, c0_n373_W_in, c0_n374_W_in, c0_n375_W_in, c0_n376_W_in, c0_n377_W_in, c0_n378_W_in, c0_n379_W_in, c0_n380_W_in, c0_n381_W_in, c0_n382_W_in, c0_n383_W_in, c0_n384_W_in, c0_n385_W_in, c0_n386_W_in, c0_n387_W_in, c0_n388_W_in, c0_n389_W_in, c0_n390_W_in, c0_n391_W_in, c0_n392_W_in, c0_n393_W_in, c0_n394_W_in, c0_n395_W_in, c0_n396_W_in, c0_n397_W_in, c0_n398_W_in, c0_n399_W_in, c0_n400_W_in, c0_n401_W_in, c0_n402_W_in, c0_n403_W_in, c0_n404_W_in, c0_n405_W_in, c0_n406_W_in, c0_n407_W_in, c0_n408_W_in, c0_n409_W_in, c0_n410_W_in, c0_n411_W_in, c0_n412_W_in, c0_n413_W_in, c0_n414_W_in, c0_n415_W_in, c0_n416_W_in, c0_n417_W_in, c0_n418_W_in, c0_n419_W_in, c0_n420_W_in, c0_n421_W_in, c0_n422_W_in, c0_n423_W_in, c0_n424_W_in, c0_n425_W_in, c0_n426_W_in, c0_n427_W_in, c0_n428_W_in, c0_n429_W_in, c0_n430_W_in, c0_n431_W_in, c0_n432_W_in, c0_n433_W_in, c0_n434_W_in, c0_n435_W_in, c0_n436_W_in, c0_n437_W_in, c0_n438_W_in, c0_n439_W_in, c0_n440_W_in, c0_n441_W_in, c0_n442_W_in, c0_n443_W_in, c0_n444_W_in, c0_n445_W_in, c0_n446_W_in, c0_n447_W_in, c0_n448_W_in, c0_n449_W_in, c0_n450_W_in, c0_n451_W_in, c0_n452_W_in, c0_n453_W_in, c0_n454_W_in, c0_n455_W_in, c0_n456_W_in, c0_n457_W_in, c0_n458_W_in, c0_n459_W_in, c0_n460_W_in, c0_n461_W_in, c0_n462_W_in, c0_n463_W_in, c0_n464_W_in, c0_n465_W_in, c0_n466_W_in, c0_n467_W_in, c0_n468_W_in, c0_n469_W_in, c0_n470_W_in, c0_n471_W_in, c0_n472_W_in, c0_n473_W_in, c0_n474_W_in, c0_n475_W_in, c0_n476_W_in, c0_n477_W_in, c0_n478_W_in, c0_n479_W_in, c0_n480_W_in, c0_n481_W_in, c0_n482_W_in, c0_n483_W_in, c0_n484_W_in, c0_n485_W_in, c0_n486_W_in, c0_n487_W_in, c0_n488_W_in, c0_n489_W_in, c0_n490_W_in, c0_n491_W_in, c0_n492_W_in, c0_n493_W_in, c0_n494_W_in, c0_n495_W_in, c0_n496_W_in, c0_n497_W_in, c0_n498_W_in, c0_n499_W_in: IN signed(BITS - 1 DOWNTO 0);
      ----------------------------------------------
      c4_n0_IO_out, c4_n1_IO_out, c4_n2_IO_out, c4_n3_IO_out, c4_n4_IO_out, c4_n5_IO_out, c4_n6_IO_out, c4_n7_IO_out, c4_n8_IO_out, c4_n9_IO_out, c4_n10_IO_out, c4_n11_IO_out, c4_n12_IO_out, c4_n13_IO_out, c4_n14_IO_out, c4_n15_IO_out, c4_n16_IO_out, c4_n17_IO_out, c4_n18_IO_out, c4_n19_IO_out, c4_n20_IO_out, c4_n21_IO_out, c4_n22_IO_out, c4_n23_IO_out, c4_n24_IO_out, c4_n25_IO_out, c4_n26_IO_out, c4_n27_IO_out, c4_n28_IO_out, c4_n29_IO_out, c4_n30_IO_out, c4_n31_IO_out, c4_n32_IO_out, c4_n33_IO_out, c4_n34_IO_out, c4_n35_IO_out, c4_n36_IO_out, c4_n37_IO_out, c4_n38_IO_out, c4_n39_IO_out, c4_n40_IO_out, c4_n41_IO_out, c4_n42_IO_out, c4_n43_IO_out, c4_n44_IO_out, c4_n45_IO_out, c4_n46_IO_out, c4_n47_IO_out, c4_n48_IO_out, c4_n49_IO_out, c4_n50_IO_out, c4_n51_IO_out, c4_n52_IO_out, c4_n53_IO_out, c4_n54_IO_out, c4_n55_IO_out, c4_n56_IO_out, c4_n57_IO_out, c4_n58_IO_out, c4_n59_IO_out, c4_n60_IO_out, c4_n61_IO_out, c4_n62_IO_out, c4_n63_IO_out, c4_n64_IO_out, c4_n65_IO_out, c4_n66_IO_out, c4_n67_IO_out, c4_n68_IO_out, c4_n69_IO_out, c4_n70_IO_out, c4_n71_IO_out, c4_n72_IO_out, c4_n73_IO_out, c4_n74_IO_out, c4_n75_IO_out, c4_n76_IO_out, c4_n77_IO_out, c4_n78_IO_out, c4_n79_IO_out, c4_n80_IO_out, c4_n81_IO_out, c4_n82_IO_out, c4_n83_IO_out, c4_n84_IO_out, c4_n85_IO_out, c4_n86_IO_out, c4_n87_IO_out, c4_n88_IO_out, c4_n89_IO_out, c4_n90_IO_out, c4_n91_IO_out, c4_n92_IO_out, c4_n93_IO_out, c4_n94_IO_out, c4_n95_IO_out, c4_n96_IO_out, c4_n97_IO_out, c4_n98_IO_out, c4_n99_IO_out, c4_n100_IO_out, c4_n101_IO_out, c4_n102_IO_out, c4_n103_IO_out, c4_n104_IO_out, c4_n105_IO_out, c4_n106_IO_out, c4_n107_IO_out, c4_n108_IO_out, c4_n109_IO_out, c4_n110_IO_out, c4_n111_IO_out, c4_n112_IO_out, c4_n113_IO_out, c4_n114_IO_out, c4_n115_IO_out, c4_n116_IO_out, c4_n117_IO_out, c4_n118_IO_out, c4_n119_IO_out, c4_n120_IO_out, c4_n121_IO_out, c4_n122_IO_out, c4_n123_IO_out, c4_n124_IO_out, c4_n125_IO_out, c4_n126_IO_out, c4_n127_IO_out, c4_n128_IO_out, c4_n129_IO_out, c4_n130_IO_out, c4_n131_IO_out, c4_n132_IO_out, c4_n133_IO_out, c4_n134_IO_out, c4_n135_IO_out, c4_n136_IO_out, c4_n137_IO_out, c4_n138_IO_out, c4_n139_IO_out, c4_n140_IO_out, c4_n141_IO_out, c4_n142_IO_out, c4_n143_IO_out, c4_n144_IO_out, c4_n145_IO_out, c4_n146_IO_out, c4_n147_IO_out, c4_n148_IO_out, c4_n149_IO_out, c4_n150_IO_out, c4_n151_IO_out, c4_n152_IO_out, c4_n153_IO_out, c4_n154_IO_out, c4_n155_IO_out, c4_n156_IO_out, c4_n157_IO_out, c4_n158_IO_out, c4_n159_IO_out, c4_n160_IO_out, c4_n161_IO_out, c4_n162_IO_out, c4_n163_IO_out, c4_n164_IO_out, c4_n165_IO_out, c4_n166_IO_out, c4_n167_IO_out, c4_n168_IO_out, c4_n169_IO_out, c4_n170_IO_out, c4_n171_IO_out, c4_n172_IO_out, c4_n173_IO_out, c4_n174_IO_out, c4_n175_IO_out, c4_n176_IO_out, c4_n177_IO_out, c4_n178_IO_out, c4_n179_IO_out, c4_n180_IO_out, c4_n181_IO_out, c4_n182_IO_out, c4_n183_IO_out, c4_n184_IO_out, c4_n185_IO_out, c4_n186_IO_out, c4_n187_IO_out, c4_n188_IO_out, c4_n189_IO_out, c4_n190_IO_out, c4_n191_IO_out, c4_n192_IO_out, c4_n193_IO_out, c4_n194_IO_out, c4_n195_IO_out, c4_n196_IO_out, c4_n197_IO_out, c4_n198_IO_out, c4_n199_IO_out, c4_n200_IO_out, c4_n201_IO_out, c4_n202_IO_out, c4_n203_IO_out, c4_n204_IO_out, c4_n205_IO_out, c4_n206_IO_out, c4_n207_IO_out, c4_n208_IO_out, c4_n209_IO_out, c4_n210_IO_out, c4_n211_IO_out, c4_n212_IO_out, c4_n213_IO_out, c4_n214_IO_out, c4_n215_IO_out, c4_n216_IO_out, c4_n217_IO_out, c4_n218_IO_out, c4_n219_IO_out, c4_n220_IO_out, c4_n221_IO_out, c4_n222_IO_out, c4_n223_IO_out, c4_n224_IO_out, c4_n225_IO_out, c4_n226_IO_out, c4_n227_IO_out, c4_n228_IO_out, c4_n229_IO_out, c4_n230_IO_out, c4_n231_IO_out, c4_n232_IO_out, c4_n233_IO_out, c4_n234_IO_out, c4_n235_IO_out, c4_n236_IO_out, c4_n237_IO_out, c4_n238_IO_out, c4_n239_IO_out, c4_n240_IO_out, c4_n241_IO_out, c4_n242_IO_out, c4_n243_IO_out, c4_n244_IO_out, c4_n245_IO_out, c4_n246_IO_out, c4_n247_IO_out, c4_n248_IO_out, c4_n249_IO_out, c4_n250_IO_out, c4_n251_IO_out, c4_n252_IO_out, c4_n253_IO_out, c4_n254_IO_out, c4_n255_IO_out, c4_n256_IO_out, c4_n257_IO_out, c4_n258_IO_out, c4_n259_IO_out, c4_n260_IO_out, c4_n261_IO_out, c4_n262_IO_out, c4_n263_IO_out, c4_n264_IO_out, c4_n265_IO_out, c4_n266_IO_out, c4_n267_IO_out, c4_n268_IO_out, c4_n269_IO_out, c4_n270_IO_out, c4_n271_IO_out, c4_n272_IO_out, c4_n273_IO_out, c4_n274_IO_out, c4_n275_IO_out, c4_n276_IO_out, c4_n277_IO_out, c4_n278_IO_out, c4_n279_IO_out, c4_n280_IO_out, c4_n281_IO_out, c4_n282_IO_out, c4_n283_IO_out, c4_n284_IO_out, c4_n285_IO_out, c4_n286_IO_out, c4_n287_IO_out, c4_n288_IO_out, c4_n289_IO_out, c4_n290_IO_out, c4_n291_IO_out, c4_n292_IO_out, c4_n293_IO_out, c4_n294_IO_out, c4_n295_IO_out, c4_n296_IO_out, c4_n297_IO_out, c4_n298_IO_out, c4_n299_IO_out, c4_n300_IO_out, c4_n301_IO_out, c4_n302_IO_out, c4_n303_IO_out, c4_n304_IO_out, c4_n305_IO_out, c4_n306_IO_out, c4_n307_IO_out, c4_n308_IO_out, c4_n309_IO_out, c4_n310_IO_out, c4_n311_IO_out, c4_n312_IO_out, c4_n313_IO_out, c4_n314_IO_out, c4_n315_IO_out, c4_n316_IO_out, c4_n317_IO_out, c4_n318_IO_out, c4_n319_IO_out, c4_n320_IO_out, c4_n321_IO_out, c4_n322_IO_out, c4_n323_IO_out, c4_n324_IO_out, c4_n325_IO_out, c4_n326_IO_out, c4_n327_IO_out, c4_n328_IO_out, c4_n329_IO_out, c4_n330_IO_out, c4_n331_IO_out, c4_n332_IO_out, c4_n333_IO_out, c4_n334_IO_out, c4_n335_IO_out, c4_n336_IO_out, c4_n337_IO_out, c4_n338_IO_out, c4_n339_IO_out, c4_n340_IO_out, c4_n341_IO_out, c4_n342_IO_out, c4_n343_IO_out, c4_n344_IO_out, c4_n345_IO_out, c4_n346_IO_out, c4_n347_IO_out, c4_n348_IO_out, c4_n349_IO_out, c4_n350_IO_out, c4_n351_IO_out, c4_n352_IO_out, c4_n353_IO_out, c4_n354_IO_out, c4_n355_IO_out, c4_n356_IO_out, c4_n357_IO_out, c4_n358_IO_out, c4_n359_IO_out, c4_n360_IO_out, c4_n361_IO_out, c4_n362_IO_out, c4_n363_IO_out, c4_n364_IO_out, c4_n365_IO_out, c4_n366_IO_out, c4_n367_IO_out, c4_n368_IO_out, c4_n369_IO_out, c4_n370_IO_out, c4_n371_IO_out, c4_n372_IO_out, c4_n373_IO_out, c4_n374_IO_out, c4_n375_IO_out, c4_n376_IO_out, c4_n377_IO_out, c4_n378_IO_out, c4_n379_IO_out, c4_n380_IO_out, c4_n381_IO_out, c4_n382_IO_out, c4_n383_IO_out, c4_n384_IO_out, c4_n385_IO_out, c4_n386_IO_out, c4_n387_IO_out, c4_n388_IO_out, c4_n389_IO_out, c4_n390_IO_out, c4_n391_IO_out, c4_n392_IO_out, c4_n393_IO_out, c4_n394_IO_out, c4_n395_IO_out, c4_n396_IO_out, c4_n397_IO_out, c4_n398_IO_out, c4_n399_IO_out, c4_n400_IO_out, c4_n401_IO_out, c4_n402_IO_out, c4_n403_IO_out, c4_n404_IO_out, c4_n405_IO_out, c4_n406_IO_out, c4_n407_IO_out, c4_n408_IO_out, c4_n409_IO_out, c4_n410_IO_out, c4_n411_IO_out, c4_n412_IO_out, c4_n413_IO_out, c4_n414_IO_out, c4_n415_IO_out, c4_n416_IO_out, c4_n417_IO_out, c4_n418_IO_out, c4_n419_IO_out, c4_n420_IO_out, c4_n421_IO_out, c4_n422_IO_out, c4_n423_IO_out, c4_n424_IO_out, c4_n425_IO_out, c4_n426_IO_out, c4_n427_IO_out, c4_n428_IO_out, c4_n429_IO_out, c4_n430_IO_out, c4_n431_IO_out, c4_n432_IO_out, c4_n433_IO_out, c4_n434_IO_out, c4_n435_IO_out, c4_n436_IO_out, c4_n437_IO_out, c4_n438_IO_out, c4_n439_IO_out, c4_n440_IO_out, c4_n441_IO_out, c4_n442_IO_out, c4_n443_IO_out, c4_n444_IO_out, c4_n445_IO_out, c4_n446_IO_out, c4_n447_IO_out, c4_n448_IO_out, c4_n449_IO_out, c4_n450_IO_out, c4_n451_IO_out, c4_n452_IO_out, c4_n453_IO_out, c4_n454_IO_out, c4_n455_IO_out, c4_n456_IO_out, c4_n457_IO_out, c4_n458_IO_out, c4_n459_IO_out, c4_n460_IO_out, c4_n461_IO_out, c4_n462_IO_out, c4_n463_IO_out, c4_n464_IO_out, c4_n465_IO_out, c4_n466_IO_out, c4_n467_IO_out, c4_n468_IO_out, c4_n469_IO_out, c4_n470_IO_out, c4_n471_IO_out, c4_n472_IO_out, c4_n473_IO_out, c4_n474_IO_out, c4_n475_IO_out, c4_n476_IO_out, c4_n477_IO_out, c4_n478_IO_out, c4_n479_IO_out, c4_n480_IO_out, c4_n481_IO_out, c4_n482_IO_out, c4_n483_IO_out, c4_n484_IO_out, c4_n485_IO_out, c4_n486_IO_out, c4_n487_IO_out, c4_n488_IO_out, c4_n489_IO_out, c4_n490_IO_out, c4_n491_IO_out, c4_n492_IO_out, c4_n493_IO_out, c4_n494_IO_out, c4_n495_IO_out, c4_n496_IO_out, c4_n497_IO_out, c4_n498_IO_out, c4_n499_IO_out: OUT signed(7 DOWNTO 0)
  );
  end ENTITY;

ARCHITECTURE arch OF  top  IS
-- SIGNALS
  SIGNAL c0_n0_W_out, c0_n1_W_out, c0_n2_W_out, c0_n3_W_out, c0_n4_W_out, c0_n5_W_out, c0_n6_W_out, c0_n7_W_out, c0_n8_W_out, c0_n9_W_out, c0_n10_W_out, c0_n11_W_out, c0_n12_W_out, c0_n13_W_out, c0_n14_W_out, c0_n15_W_out, c0_n16_W_out, c0_n17_W_out, c0_n18_W_out, c0_n19_W_out, c0_n20_W_out, c0_n21_W_out, c0_n22_W_out, c0_n23_W_out, c0_n24_W_out, c0_n25_W_out, c0_n26_W_out, c0_n27_W_out, c0_n28_W_out, c0_n29_W_out, c0_n30_W_out, c0_n31_W_out, c0_n32_W_out, c0_n33_W_out, c0_n34_W_out, c0_n35_W_out, c0_n36_W_out, c0_n37_W_out, c0_n38_W_out, c0_n39_W_out, c0_n40_W_out, c0_n41_W_out, c0_n42_W_out, c0_n43_W_out, c0_n44_W_out, c0_n45_W_out, c0_n46_W_out, c0_n47_W_out, c0_n48_W_out, c0_n49_W_out, c0_n50_W_out, c0_n51_W_out, c0_n52_W_out, c0_n53_W_out, c0_n54_W_out, c0_n55_W_out, c0_n56_W_out, c0_n57_W_out, c0_n58_W_out, c0_n59_W_out, c0_n60_W_out, c0_n61_W_out, c0_n62_W_out, c0_n63_W_out, c0_n64_W_out, c0_n65_W_out, c0_n66_W_out, c0_n67_W_out, c0_n68_W_out, c0_n69_W_out, c0_n70_W_out, c0_n71_W_out, c0_n72_W_out, c0_n73_W_out, c0_n74_W_out, c0_n75_W_out, c0_n76_W_out, c0_n77_W_out, c0_n78_W_out, c0_n79_W_out, c0_n80_W_out, c0_n81_W_out, c0_n82_W_out, c0_n83_W_out, c0_n84_W_out, c0_n85_W_out, c0_n86_W_out, c0_n87_W_out, c0_n88_W_out, c0_n89_W_out, c0_n90_W_out, c0_n91_W_out, c0_n92_W_out, c0_n93_W_out, c0_n94_W_out, c0_n95_W_out, c0_n96_W_out, c0_n97_W_out, c0_n98_W_out, c0_n99_W_out, c0_n100_W_out, c0_n101_W_out, c0_n102_W_out, c0_n103_W_out, c0_n104_W_out, c0_n105_W_out, c0_n106_W_out, c0_n107_W_out, c0_n108_W_out, c0_n109_W_out, c0_n110_W_out, c0_n111_W_out, c0_n112_W_out, c0_n113_W_out, c0_n114_W_out, c0_n115_W_out, c0_n116_W_out, c0_n117_W_out, c0_n118_W_out, c0_n119_W_out, c0_n120_W_out, c0_n121_W_out, c0_n122_W_out, c0_n123_W_out, c0_n124_W_out, c0_n125_W_out, c0_n126_W_out, c0_n127_W_out, c0_n128_W_out, c0_n129_W_out, c0_n130_W_out, c0_n131_W_out, c0_n132_W_out, c0_n133_W_out, c0_n134_W_out, c0_n135_W_out, c0_n136_W_out, c0_n137_W_out, c0_n138_W_out, c0_n139_W_out, c0_n140_W_out, c0_n141_W_out, c0_n142_W_out, c0_n143_W_out, c0_n144_W_out, c0_n145_W_out, c0_n146_W_out, c0_n147_W_out, c0_n148_W_out, c0_n149_W_out, c0_n150_W_out, c0_n151_W_out, c0_n152_W_out, c0_n153_W_out, c0_n154_W_out, c0_n155_W_out, c0_n156_W_out, c0_n157_W_out, c0_n158_W_out, c0_n159_W_out, c0_n160_W_out, c0_n161_W_out, c0_n162_W_out, c0_n163_W_out, c0_n164_W_out, c0_n165_W_out, c0_n166_W_out, c0_n167_W_out, c0_n168_W_out, c0_n169_W_out, c0_n170_W_out, c0_n171_W_out, c0_n172_W_out, c0_n173_W_out, c0_n174_W_out, c0_n175_W_out, c0_n176_W_out, c0_n177_W_out, c0_n178_W_out, c0_n179_W_out, c0_n180_W_out, c0_n181_W_out, c0_n182_W_out, c0_n183_W_out, c0_n184_W_out, c0_n185_W_out, c0_n186_W_out, c0_n187_W_out, c0_n188_W_out, c0_n189_W_out, c0_n190_W_out, c0_n191_W_out, c0_n192_W_out, c0_n193_W_out, c0_n194_W_out, c0_n195_W_out, c0_n196_W_out, c0_n197_W_out, c0_n198_W_out, c0_n199_W_out, c0_n200_W_out, c0_n201_W_out, c0_n202_W_out, c0_n203_W_out, c0_n204_W_out, c0_n205_W_out, c0_n206_W_out, c0_n207_W_out, c0_n208_W_out, c0_n209_W_out, c0_n210_W_out, c0_n211_W_out, c0_n212_W_out, c0_n213_W_out, c0_n214_W_out, c0_n215_W_out, c0_n216_W_out, c0_n217_W_out, c0_n218_W_out, c0_n219_W_out, c0_n220_W_out, c0_n221_W_out, c0_n222_W_out, c0_n223_W_out, c0_n224_W_out, c0_n225_W_out, c0_n226_W_out, c0_n227_W_out, c0_n228_W_out, c0_n229_W_out, c0_n230_W_out, c0_n231_W_out, c0_n232_W_out, c0_n233_W_out, c0_n234_W_out, c0_n235_W_out, c0_n236_W_out, c0_n237_W_out, c0_n238_W_out, c0_n239_W_out, c0_n240_W_out, c0_n241_W_out, c0_n242_W_out, c0_n243_W_out, c0_n244_W_out, c0_n245_W_out, c0_n246_W_out, c0_n247_W_out, c0_n248_W_out, c0_n249_W_out, c0_n250_W_out, c0_n251_W_out, c0_n252_W_out, c0_n253_W_out, c0_n254_W_out, c0_n255_W_out, c0_n256_W_out, c0_n257_W_out, c0_n258_W_out, c0_n259_W_out, c0_n260_W_out, c0_n261_W_out, c0_n262_W_out, c0_n263_W_out, c0_n264_W_out, c0_n265_W_out, c0_n266_W_out, c0_n267_W_out, c0_n268_W_out, c0_n269_W_out, c0_n270_W_out, c0_n271_W_out, c0_n272_W_out, c0_n273_W_out, c0_n274_W_out, c0_n275_W_out, c0_n276_W_out, c0_n277_W_out, c0_n278_W_out, c0_n279_W_out, c0_n280_W_out, c0_n281_W_out, c0_n282_W_out, c0_n283_W_out, c0_n284_W_out, c0_n285_W_out, c0_n286_W_out, c0_n287_W_out, c0_n288_W_out, c0_n289_W_out, c0_n290_W_out, c0_n291_W_out, c0_n292_W_out, c0_n293_W_out, c0_n294_W_out, c0_n295_W_out, c0_n296_W_out, c0_n297_W_out, c0_n298_W_out, c0_n299_W_out, c0_n300_W_out, c0_n301_W_out, c0_n302_W_out, c0_n303_W_out, c0_n304_W_out, c0_n305_W_out, c0_n306_W_out, c0_n307_W_out, c0_n308_W_out, c0_n309_W_out, c0_n310_W_out, c0_n311_W_out, c0_n312_W_out, c0_n313_W_out, c0_n314_W_out, c0_n315_W_out, c0_n316_W_out, c0_n317_W_out, c0_n318_W_out, c0_n319_W_out, c0_n320_W_out, c0_n321_W_out, c0_n322_W_out, c0_n323_W_out, c0_n324_W_out, c0_n325_W_out, c0_n326_W_out, c0_n327_W_out, c0_n328_W_out, c0_n329_W_out, c0_n330_W_out, c0_n331_W_out, c0_n332_W_out, c0_n333_W_out, c0_n334_W_out, c0_n335_W_out, c0_n336_W_out, c0_n337_W_out, c0_n338_W_out, c0_n339_W_out, c0_n340_W_out, c0_n341_W_out, c0_n342_W_out, c0_n343_W_out, c0_n344_W_out, c0_n345_W_out, c0_n346_W_out, c0_n347_W_out, c0_n348_W_out, c0_n349_W_out, c0_n350_W_out, c0_n351_W_out, c0_n352_W_out, c0_n353_W_out, c0_n354_W_out, c0_n355_W_out, c0_n356_W_out, c0_n357_W_out, c0_n358_W_out, c0_n359_W_out, c0_n360_W_out, c0_n361_W_out, c0_n362_W_out, c0_n363_W_out, c0_n364_W_out, c0_n365_W_out, c0_n366_W_out, c0_n367_W_out, c0_n368_W_out, c0_n369_W_out, c0_n370_W_out, c0_n371_W_out, c0_n372_W_out, c0_n373_W_out, c0_n374_W_out, c0_n375_W_out, c0_n376_W_out, c0_n377_W_out, c0_n378_W_out, c0_n379_W_out, c0_n380_W_out, c0_n381_W_out, c0_n382_W_out, c0_n383_W_out, c0_n384_W_out, c0_n385_W_out, c0_n386_W_out, c0_n387_W_out, c0_n388_W_out, c0_n389_W_out, c0_n390_W_out, c0_n391_W_out, c0_n392_W_out, c0_n393_W_out, c0_n394_W_out, c0_n395_W_out, c0_n396_W_out, c0_n397_W_out, c0_n398_W_out, c0_n399_W_out, c0_n400_W_out, c0_n401_W_out, c0_n402_W_out, c0_n403_W_out, c0_n404_W_out, c0_n405_W_out, c0_n406_W_out, c0_n407_W_out, c0_n408_W_out, c0_n409_W_out, c0_n410_W_out, c0_n411_W_out, c0_n412_W_out, c0_n413_W_out, c0_n414_W_out, c0_n415_W_out, c0_n416_W_out, c0_n417_W_out, c0_n418_W_out, c0_n419_W_out, c0_n420_W_out, c0_n421_W_out, c0_n422_W_out, c0_n423_W_out, c0_n424_W_out, c0_n425_W_out, c0_n426_W_out, c0_n427_W_out, c0_n428_W_out, c0_n429_W_out, c0_n430_W_out, c0_n431_W_out, c0_n432_W_out, c0_n433_W_out, c0_n434_W_out, c0_n435_W_out, c0_n436_W_out, c0_n437_W_out, c0_n438_W_out, c0_n439_W_out, c0_n440_W_out, c0_n441_W_out, c0_n442_W_out, c0_n443_W_out, c0_n444_W_out, c0_n445_W_out, c0_n446_W_out, c0_n447_W_out, c0_n448_W_out, c0_n449_W_out, c0_n450_W_out, c0_n451_W_out, c0_n452_W_out, c0_n453_W_out, c0_n454_W_out, c0_n455_W_out, c0_n456_W_out, c0_n457_W_out, c0_n458_W_out, c0_n459_W_out, c0_n460_W_out, c0_n461_W_out, c0_n462_W_out, c0_n463_W_out, c0_n464_W_out, c0_n465_W_out, c0_n466_W_out, c0_n467_W_out, c0_n468_W_out, c0_n469_W_out, c0_n470_W_out, c0_n471_W_out, c0_n472_W_out, c0_n473_W_out, c0_n474_W_out, c0_n475_W_out, c0_n476_W_out, c0_n477_W_out, c0_n478_W_out, c0_n479_W_out, c0_n480_W_out, c0_n481_W_out, c0_n482_W_out, c0_n483_W_out, c0_n484_W_out, c0_n485_W_out, c0_n486_W_out, c0_n487_W_out, c0_n488_W_out, c0_n489_W_out, c0_n490_W_out, c0_n491_W_out, c0_n492_W_out, c0_n493_W_out, c0_n494_W_out, c0_n495_W_out, c0_n496_W_out, c0_n497_W_out, c0_n498_W_out, c0_n499_W_out, c1_n0_W_out, c1_n1_W_out, c1_n2_W_out, c1_n3_W_out, c1_n4_W_out, c1_n5_W_out, c1_n6_W_out, c1_n7_W_out, c1_n8_W_out, c1_n9_W_out, c1_n10_W_out, c1_n11_W_out, c1_n12_W_out, c1_n13_W_out, c1_n14_W_out, c1_n15_W_out, c1_n16_W_out, c1_n17_W_out, c1_n18_W_out, c1_n19_W_out, c1_n20_W_out, c1_n21_W_out, c1_n22_W_out, c1_n23_W_out, c1_n24_W_out, c1_n25_W_out, c1_n26_W_out, c1_n27_W_out, c1_n28_W_out, c1_n29_W_out, c1_n30_W_out, c1_n31_W_out, c1_n32_W_out, c1_n33_W_out, c1_n34_W_out, c1_n35_W_out, c1_n36_W_out, c1_n37_W_out, c1_n38_W_out, c1_n39_W_out, c1_n40_W_out, c1_n41_W_out, c1_n42_W_out, c1_n43_W_out, c1_n44_W_out, c1_n45_W_out, c1_n46_W_out, c1_n47_W_out, c1_n48_W_out, c1_n49_W_out, c1_n50_W_out, c1_n51_W_out, c1_n52_W_out, c1_n53_W_out, c1_n54_W_out, c1_n55_W_out, c1_n56_W_out, c1_n57_W_out, c1_n58_W_out, c1_n59_W_out, c1_n60_W_out, c1_n61_W_out, c1_n62_W_out, c1_n63_W_out, c1_n64_W_out, c1_n65_W_out, c1_n66_W_out, c1_n67_W_out, c1_n68_W_out, c1_n69_W_out, c1_n70_W_out, c1_n71_W_out, c1_n72_W_out, c1_n73_W_out, c1_n74_W_out, c1_n75_W_out, c1_n76_W_out, c1_n77_W_out, c1_n78_W_out, c1_n79_W_out, c1_n80_W_out, c1_n81_W_out, c1_n82_W_out, c1_n83_W_out, c1_n84_W_out, c1_n85_W_out, c1_n86_W_out, c1_n87_W_out, c1_n88_W_out, c1_n89_W_out, c1_n90_W_out, c1_n91_W_out, c1_n92_W_out, c1_n93_W_out, c1_n94_W_out, c1_n95_W_out, c1_n96_W_out, c1_n97_W_out, c1_n98_W_out, c1_n99_W_out, c1_n100_W_out, c1_n101_W_out, c1_n102_W_out, c1_n103_W_out, c1_n104_W_out, c1_n105_W_out, c1_n106_W_out, c1_n107_W_out, c1_n108_W_out, c1_n109_W_out, c1_n110_W_out, c1_n111_W_out, c1_n112_W_out, c1_n113_W_out, c1_n114_W_out, c1_n115_W_out, c1_n116_W_out, c1_n117_W_out, c1_n118_W_out, c1_n119_W_out, c1_n120_W_out, c1_n121_W_out, c1_n122_W_out, c1_n123_W_out, c1_n124_W_out, c1_n125_W_out, c1_n126_W_out, c1_n127_W_out, c1_n128_W_out, c1_n129_W_out, c1_n130_W_out, c1_n131_W_out, c1_n132_W_out, c1_n133_W_out, c1_n134_W_out, c1_n135_W_out, c1_n136_W_out, c1_n137_W_out, c1_n138_W_out, c1_n139_W_out, c1_n140_W_out, c1_n141_W_out, c1_n142_W_out, c1_n143_W_out, c1_n144_W_out, c1_n145_W_out, c1_n146_W_out, c1_n147_W_out, c1_n148_W_out, c1_n149_W_out, c1_n150_W_out, c1_n151_W_out, c1_n152_W_out, c1_n153_W_out, c1_n154_W_out, c1_n155_W_out, c1_n156_W_out, c1_n157_W_out, c1_n158_W_out, c1_n159_W_out, c1_n160_W_out, c1_n161_W_out, c1_n162_W_out, c1_n163_W_out, c1_n164_W_out, c1_n165_W_out, c1_n166_W_out, c1_n167_W_out, c1_n168_W_out, c1_n169_W_out, c1_n170_W_out, c1_n171_W_out, c1_n172_W_out, c1_n173_W_out, c1_n174_W_out, c1_n175_W_out, c1_n176_W_out, c1_n177_W_out, c1_n178_W_out, c1_n179_W_out, c1_n180_W_out, c1_n181_W_out, c1_n182_W_out, c1_n183_W_out, c1_n184_W_out, c1_n185_W_out, c1_n186_W_out, c1_n187_W_out, c1_n188_W_out, c1_n189_W_out, c1_n190_W_out, c1_n191_W_out, c1_n192_W_out, c1_n193_W_out, c1_n194_W_out, c1_n195_W_out, c1_n196_W_out, c1_n197_W_out, c1_n198_W_out, c1_n199_W_out, c1_n200_W_out, c1_n201_W_out, c1_n202_W_out, c1_n203_W_out, c1_n204_W_out, c1_n205_W_out, c1_n206_W_out, c1_n207_W_out, c1_n208_W_out, c1_n209_W_out, c1_n210_W_out, c1_n211_W_out, c1_n212_W_out, c1_n213_W_out, c1_n214_W_out, c1_n215_W_out, c1_n216_W_out, c1_n217_W_out, c1_n218_W_out, c1_n219_W_out, c1_n220_W_out, c1_n221_W_out, c1_n222_W_out, c1_n223_W_out, c1_n224_W_out, c1_n225_W_out, c1_n226_W_out, c1_n227_W_out, c1_n228_W_out, c1_n229_W_out, c1_n230_W_out, c1_n231_W_out, c1_n232_W_out, c1_n233_W_out, c1_n234_W_out, c1_n235_W_out, c1_n236_W_out, c1_n237_W_out, c1_n238_W_out, c1_n239_W_out, c1_n240_W_out, c1_n241_W_out, c1_n242_W_out, c1_n243_W_out, c1_n244_W_out, c1_n245_W_out, c1_n246_W_out, c1_n247_W_out, c1_n248_W_out, c1_n249_W_out, c1_n250_W_out, c1_n251_W_out, c1_n252_W_out, c1_n253_W_out, c1_n254_W_out, c1_n255_W_out, c1_n256_W_out, c1_n257_W_out, c1_n258_W_out, c1_n259_W_out, c1_n260_W_out, c1_n261_W_out, c1_n262_W_out, c1_n263_W_out, c1_n264_W_out, c1_n265_W_out, c1_n266_W_out, c1_n267_W_out, c1_n268_W_out, c1_n269_W_out, c1_n270_W_out, c1_n271_W_out, c1_n272_W_out, c1_n273_W_out, c1_n274_W_out, c1_n275_W_out, c1_n276_W_out, c1_n277_W_out, c1_n278_W_out, c1_n279_W_out, c1_n280_W_out, c1_n281_W_out, c1_n282_W_out, c1_n283_W_out, c1_n284_W_out, c1_n285_W_out, c1_n286_W_out, c1_n287_W_out, c1_n288_W_out, c1_n289_W_out, c1_n290_W_out, c1_n291_W_out, c1_n292_W_out, c1_n293_W_out, c1_n294_W_out, c1_n295_W_out, c1_n296_W_out, c1_n297_W_out, c1_n298_W_out, c1_n299_W_out, c2_n0_W_out, c2_n1_W_out, c2_n2_W_out, c2_n3_W_out, c2_n4_W_out, c2_n5_W_out, c2_n6_W_out, c2_n7_W_out, c2_n8_W_out, c2_n9_W_out, c2_n10_W_out, c2_n11_W_out, c2_n12_W_out, c2_n13_W_out, c2_n14_W_out, c2_n15_W_out, c2_n16_W_out, c2_n17_W_out, c2_n18_W_out, c2_n19_W_out, c2_n20_W_out, c2_n21_W_out, c2_n22_W_out, c2_n23_W_out, c2_n24_W_out, c2_n25_W_out, c2_n26_W_out, c2_n27_W_out, c2_n28_W_out, c2_n29_W_out, c2_n30_W_out, c2_n31_W_out, c2_n32_W_out, c2_n33_W_out, c2_n34_W_out, c2_n35_W_out, c2_n36_W_out, c2_n37_W_out, c2_n38_W_out, c2_n39_W_out, c2_n40_W_out, c2_n41_W_out, c2_n42_W_out, c2_n43_W_out, c2_n44_W_out, c2_n45_W_out, c2_n46_W_out, c2_n47_W_out, c2_n48_W_out, c2_n49_W_out, c2_n50_W_out, c2_n51_W_out, c2_n52_W_out, c2_n53_W_out, c2_n54_W_out, c2_n55_W_out, c2_n56_W_out, c2_n57_W_out, c2_n58_W_out, c2_n59_W_out, c2_n60_W_out, c2_n61_W_out, c2_n62_W_out, c2_n63_W_out, c2_n64_W_out, c2_n65_W_out, c2_n66_W_out, c2_n67_W_out, c2_n68_W_out, c2_n69_W_out, c2_n70_W_out, c2_n71_W_out, c2_n72_W_out, c2_n73_W_out, c2_n74_W_out, c2_n75_W_out, c2_n76_W_out, c2_n77_W_out, c2_n78_W_out, c2_n79_W_out, c2_n80_W_out, c2_n81_W_out, c2_n82_W_out, c2_n83_W_out, c2_n84_W_out, c2_n85_W_out, c2_n86_W_out, c2_n87_W_out, c2_n88_W_out, c2_n89_W_out, c2_n90_W_out, c2_n91_W_out, c2_n92_W_out, c2_n93_W_out, c2_n94_W_out, c2_n95_W_out, c2_n96_W_out, c2_n97_W_out, c2_n98_W_out, c2_n99_W_out, c3_n100_W_out, c3_n101_W_out, c3_n102_W_out, c3_n103_W_out, c3_n104_W_out, c3_n105_W_out, c3_n106_W_out, c3_n107_W_out, c3_n108_W_out, c3_n109_W_out, c3_n110_W_out, c3_n111_W_out, c3_n112_W_out, c3_n113_W_out, c3_n114_W_out, c3_n115_W_out, c3_n116_W_out, c3_n117_W_out, c3_n118_W_out, c3_n119_W_out, c3_n120_W_out, c3_n121_W_out, c3_n122_W_out, c3_n123_W_out, c3_n124_W_out, c3_n125_W_out, c3_n126_W_out, c3_n127_W_out, c3_n128_W_out, c3_n129_W_out, c3_n130_W_out, c3_n131_W_out, c3_n132_W_out, c3_n133_W_out, c3_n134_W_out, c3_n135_W_out, c3_n136_W_out, c3_n137_W_out, c3_n138_W_out, c3_n139_W_out, c3_n140_W_out, c3_n141_W_out, c3_n142_W_out, c3_n143_W_out, c3_n144_W_out, c3_n145_W_out, c3_n146_W_out, c3_n147_W_out, c3_n148_W_out, c3_n149_W_out, c3_n150_W_out, c3_n151_W_out, c3_n152_W_out, c3_n153_W_out, c3_n154_W_out, c3_n155_W_out, c3_n156_W_out, c3_n157_W_out, c3_n158_W_out, c3_n159_W_out, c3_n160_W_out, c3_n161_W_out, c3_n162_W_out, c3_n163_W_out, c3_n164_W_out, c3_n165_W_out, c3_n166_W_out, c3_n167_W_out, c3_n168_W_out, c3_n169_W_out, c3_n170_W_out, c3_n171_W_out, c3_n172_W_out, c3_n173_W_out, c3_n174_W_out, c3_n175_W_out, c3_n176_W_out, c3_n177_W_out, c3_n178_W_out, c3_n179_W_out, c3_n180_W_out, c3_n181_W_out, c3_n182_W_out, c3_n183_W_out, c3_n184_W_out, c3_n185_W_out, c3_n186_W_out, c3_n187_W_out, c3_n188_W_out, c3_n189_W_out, c3_n190_W_out, c3_n191_W_out, c3_n192_W_out, c3_n193_W_out, c3_n194_W_out, c3_n195_W_out, c3_n196_W_out, c3_n197_W_out, c3_n198_W_out, c3_n199_W_out, c3_n200_W_out, c3_n201_W_out, c3_n202_W_out, c3_n203_W_out, c3_n204_W_out, c3_n205_W_out, c3_n206_W_out, c3_n207_W_out, c3_n208_W_out, c3_n209_W_out, c3_n210_W_out, c3_n211_W_out, c3_n212_W_out, c3_n213_W_out, c3_n214_W_out, c3_n215_W_out, c3_n216_W_out, c3_n217_W_out, c3_n218_W_out, c3_n219_W_out, c3_n220_W_out, c3_n221_W_out, c3_n222_W_out, c3_n223_W_out, c3_n224_W_out, c3_n225_W_out, c3_n226_W_out, c3_n227_W_out, c3_n228_W_out, c3_n229_W_out, c3_n230_W_out, c3_n231_W_out, c3_n232_W_out, c3_n233_W_out, c3_n234_W_out, c3_n235_W_out, c3_n236_W_out, c3_n237_W_out, c3_n238_W_out, c3_n239_W_out, c3_n240_W_out, c3_n241_W_out, c3_n242_W_out, c3_n243_W_out, c3_n244_W_out, c3_n245_W_out, c3_n246_W_out, c3_n247_W_out, c3_n248_W_out, c3_n249_W_out, c3_n250_W_out, c3_n251_W_out, c3_n252_W_out, c3_n253_W_out, c3_n254_W_out, c3_n255_W_out, c3_n256_W_out, c3_n257_W_out, c3_n258_W_out, c3_n259_W_out, c3_n260_W_out, c3_n261_W_out, c3_n262_W_out, c3_n263_W_out, c3_n264_W_out, c3_n265_W_out, c3_n266_W_out, c3_n267_W_out, c3_n268_W_out, c3_n269_W_out, c3_n270_W_out, c3_n271_W_out, c3_n272_W_out, c3_n273_W_out, c3_n274_W_out, c3_n275_W_out, c3_n276_W_out, c3_n277_W_out, c3_n278_W_out, c3_n279_W_out, c3_n280_W_out, c3_n281_W_out, c3_n282_W_out, c3_n283_W_out, c3_n284_W_out, c3_n285_W_out, c3_n286_W_out, c3_n287_W_out, c3_n288_W_out, c3_n289_W_out, c3_n290_W_out, c3_n291_W_out, c3_n292_W_out, c3_n293_W_out, c3_n294_W_out, c3_n295_W_out, c3_n296_W_out, c3_n297_W_out, c3_n298_W_out, c3_n299_W_out, c3_n0_W_out, c3_n1_W_out, c3_n2_W_out, c3_n3_W_out, c3_n4_W_out, c3_n5_W_out, c3_n6_W_out, c3_n7_W_out, c3_n8_W_out, c3_n9_W_out, c3_n10_W_out, c3_n11_W_out, c3_n12_W_out, c3_n13_W_out, c3_n14_W_out, c3_n15_W_out, c3_n16_W_out, c3_n17_W_out, c3_n18_W_out, c3_n19_W_out, c3_n20_W_out, c3_n21_W_out, c3_n22_W_out, c3_n23_W_out, c3_n24_W_out, c3_n25_W_out, c3_n26_W_out, c3_n27_W_out, c3_n28_W_out, c3_n29_W_out, c3_n30_W_out, c3_n31_W_out, c3_n32_W_out, c3_n33_W_out, c3_n34_W_out, c3_n35_W_out, c3_n36_W_out, c3_n37_W_out, c3_n38_W_out, c3_n39_W_out, c3_n40_W_out, c3_n41_W_out, c3_n42_W_out, c3_n43_W_out, c3_n44_W_out, c3_n45_W_out, c3_n46_W_out, c3_n47_W_out, c3_n48_W_out, c3_n49_W_out, c3_n50_W_out, c3_n51_W_out, c3_n52_W_out, c3_n53_W_out, c3_n54_W_out, c3_n55_W_out, c3_n56_W_out, c3_n57_W_out, c3_n58_W_out, c3_n59_W_out, c3_n60_W_out, c3_n61_W_out, c3_n62_W_out, c3_n63_W_out, c3_n64_W_out, c3_n65_W_out, c3_n66_W_out, c3_n67_W_out, c3_n68_W_out, c3_n69_W_out, c3_n70_W_out, c3_n71_W_out, c3_n72_W_out, c3_n73_W_out, c3_n74_W_out, c3_n75_W_out, c3_n76_W_out, c3_n77_W_out, c3_n78_W_out, c3_n79_W_out, c3_n80_W_out, c3_n81_W_out, c3_n82_W_out, c3_n83_W_out, c3_n84_W_out, c3_n85_W_out, c3_n86_W_out, c3_n87_W_out, c3_n88_W_out, c3_n89_W_out, c3_n90_W_out, c3_n91_W_out, c3_n92_W_out, c3_n93_W_out, c3_n94_W_out, c3_n95_W_out, c3_n96_W_out, c3_n97_W_out, c3_n98_W_out, c3_n99_W_out: signed(BITS - 1 DOWNTO 0);
  SIGNAL c1_IO_in:  signed((BITS*500) - 1 DOWNTO 0);
  SIGNAL c2_IO_in:  signed((BITS*300) - 1 DOWNTO 0);
  SIGNAL c3_IO_in:  signed((BITS*100) - 1 DOWNTO 0);
  SIGNAL c4_IO_in:  signed((BITS*300) - 1 DOWNTO 0);
  SIGNAL c0_n0_IO_out, c0_n1_IO_out, c0_n2_IO_out, c0_n3_IO_out, c0_n4_IO_out, c0_n5_IO_out, c0_n6_IO_out, c0_n7_IO_out, c0_n8_IO_out, c0_n9_IO_out, c0_n10_IO_out, c0_n11_IO_out, c0_n12_IO_out, c0_n13_IO_out, c0_n14_IO_out, c0_n15_IO_out, c0_n16_IO_out, c0_n17_IO_out, c0_n18_IO_out, c0_n19_IO_out, c0_n20_IO_out, c0_n21_IO_out, c0_n22_IO_out, c0_n23_IO_out, c0_n24_IO_out, c0_n25_IO_out, c0_n26_IO_out, c0_n27_IO_out, c0_n28_IO_out, c0_n29_IO_out, c0_n30_IO_out, c0_n31_IO_out, c0_n32_IO_out, c0_n33_IO_out, c0_n34_IO_out, c0_n35_IO_out, c0_n36_IO_out, c0_n37_IO_out, c0_n38_IO_out, c0_n39_IO_out, c0_n40_IO_out, c0_n41_IO_out, c0_n42_IO_out, c0_n43_IO_out, c0_n44_IO_out, c0_n45_IO_out, c0_n46_IO_out, c0_n47_IO_out, c0_n48_IO_out, c0_n49_IO_out, c0_n50_IO_out, c0_n51_IO_out, c0_n52_IO_out, c0_n53_IO_out, c0_n54_IO_out, c0_n55_IO_out, c0_n56_IO_out, c0_n57_IO_out, c0_n58_IO_out, c0_n59_IO_out, c0_n60_IO_out, c0_n61_IO_out, c0_n62_IO_out, c0_n63_IO_out, c0_n64_IO_out, c0_n65_IO_out, c0_n66_IO_out, c0_n67_IO_out, c0_n68_IO_out, c0_n69_IO_out, c0_n70_IO_out, c0_n71_IO_out, c0_n72_IO_out, c0_n73_IO_out, c0_n74_IO_out, c0_n75_IO_out, c0_n76_IO_out, c0_n77_IO_out, c0_n78_IO_out, c0_n79_IO_out, c0_n80_IO_out, c0_n81_IO_out, c0_n82_IO_out, c0_n83_IO_out, c0_n84_IO_out, c0_n85_IO_out, c0_n86_IO_out, c0_n87_IO_out, c0_n88_IO_out, c0_n89_IO_out, c0_n90_IO_out, c0_n91_IO_out, c0_n92_IO_out, c0_n93_IO_out, c0_n94_IO_out, c0_n95_IO_out, c0_n96_IO_out, c0_n97_IO_out, c0_n98_IO_out, c0_n99_IO_out, c0_n100_IO_out, c0_n101_IO_out, c0_n102_IO_out, c0_n103_IO_out, c0_n104_IO_out, c0_n105_IO_out, c0_n106_IO_out, c0_n107_IO_out, c0_n108_IO_out, c0_n109_IO_out, c0_n110_IO_out, c0_n111_IO_out, c0_n112_IO_out, c0_n113_IO_out, c0_n114_IO_out, c0_n115_IO_out, c0_n116_IO_out, c0_n117_IO_out, c0_n118_IO_out, c0_n119_IO_out, c0_n120_IO_out, c0_n121_IO_out, c0_n122_IO_out, c0_n123_IO_out, c0_n124_IO_out, c0_n125_IO_out, c0_n126_IO_out, c0_n127_IO_out, c0_n128_IO_out, c0_n129_IO_out, c0_n130_IO_out, c0_n131_IO_out, c0_n132_IO_out, c0_n133_IO_out, c0_n134_IO_out, c0_n135_IO_out, c0_n136_IO_out, c0_n137_IO_out, c0_n138_IO_out, c0_n139_IO_out, c0_n140_IO_out, c0_n141_IO_out, c0_n142_IO_out, c0_n143_IO_out, c0_n144_IO_out, c0_n145_IO_out, c0_n146_IO_out, c0_n147_IO_out, c0_n148_IO_out, c0_n149_IO_out, c0_n150_IO_out, c0_n151_IO_out, c0_n152_IO_out, c0_n153_IO_out, c0_n154_IO_out, c0_n155_IO_out, c0_n156_IO_out, c0_n157_IO_out, c0_n158_IO_out, c0_n159_IO_out, c0_n160_IO_out, c0_n161_IO_out, c0_n162_IO_out, c0_n163_IO_out, c0_n164_IO_out, c0_n165_IO_out, c0_n166_IO_out, c0_n167_IO_out, c0_n168_IO_out, c0_n169_IO_out, c0_n170_IO_out, c0_n171_IO_out, c0_n172_IO_out, c0_n173_IO_out, c0_n174_IO_out, c0_n175_IO_out, c0_n176_IO_out, c0_n177_IO_out, c0_n178_IO_out, c0_n179_IO_out, c0_n180_IO_out, c0_n181_IO_out, c0_n182_IO_out, c0_n183_IO_out, c0_n184_IO_out, c0_n185_IO_out, c0_n186_IO_out, c0_n187_IO_out, c0_n188_IO_out, c0_n189_IO_out, c0_n190_IO_out, c0_n191_IO_out, c0_n192_IO_out, c0_n193_IO_out, c0_n194_IO_out, c0_n195_IO_out, c0_n196_IO_out, c0_n197_IO_out, c0_n198_IO_out, c0_n199_IO_out, c0_n200_IO_out, c0_n201_IO_out, c0_n202_IO_out, c0_n203_IO_out, c0_n204_IO_out, c0_n205_IO_out, c0_n206_IO_out, c0_n207_IO_out, c0_n208_IO_out, c0_n209_IO_out, c0_n210_IO_out, c0_n211_IO_out, c0_n212_IO_out, c0_n213_IO_out, c0_n214_IO_out, c0_n215_IO_out, c0_n216_IO_out, c0_n217_IO_out, c0_n218_IO_out, c0_n219_IO_out, c0_n220_IO_out, c0_n221_IO_out, c0_n222_IO_out, c0_n223_IO_out, c0_n224_IO_out, c0_n225_IO_out, c0_n226_IO_out, c0_n227_IO_out, c0_n228_IO_out, c0_n229_IO_out, c0_n230_IO_out, c0_n231_IO_out, c0_n232_IO_out, c0_n233_IO_out, c0_n234_IO_out, c0_n235_IO_out, c0_n236_IO_out, c0_n237_IO_out, c0_n238_IO_out, c0_n239_IO_out, c0_n240_IO_out, c0_n241_IO_out, c0_n242_IO_out, c0_n243_IO_out, c0_n244_IO_out, c0_n245_IO_out, c0_n246_IO_out, c0_n247_IO_out, c0_n248_IO_out, c0_n249_IO_out, c0_n250_IO_out, c0_n251_IO_out, c0_n252_IO_out, c0_n253_IO_out, c0_n254_IO_out, c0_n255_IO_out, c0_n256_IO_out, c0_n257_IO_out, c0_n258_IO_out, c0_n259_IO_out, c0_n260_IO_out, c0_n261_IO_out, c0_n262_IO_out, c0_n263_IO_out, c0_n264_IO_out, c0_n265_IO_out, c0_n266_IO_out, c0_n267_IO_out, c0_n268_IO_out, c0_n269_IO_out, c0_n270_IO_out, c0_n271_IO_out, c0_n272_IO_out, c0_n273_IO_out, c0_n274_IO_out, c0_n275_IO_out, c0_n276_IO_out, c0_n277_IO_out, c0_n278_IO_out, c0_n279_IO_out, c0_n280_IO_out, c0_n281_IO_out, c0_n282_IO_out, c0_n283_IO_out, c0_n284_IO_out, c0_n285_IO_out, c0_n286_IO_out, c0_n287_IO_out, c0_n288_IO_out, c0_n289_IO_out, c0_n290_IO_out, c0_n291_IO_out, c0_n292_IO_out, c0_n293_IO_out, c0_n294_IO_out, c0_n295_IO_out, c0_n296_IO_out, c0_n297_IO_out, c0_n298_IO_out, c0_n299_IO_out, c0_n300_IO_out, c0_n301_IO_out, c0_n302_IO_out, c0_n303_IO_out, c0_n304_IO_out, c0_n305_IO_out, c0_n306_IO_out, c0_n307_IO_out, c0_n308_IO_out, c0_n309_IO_out, c0_n310_IO_out, c0_n311_IO_out, c0_n312_IO_out, c0_n313_IO_out, c0_n314_IO_out, c0_n315_IO_out, c0_n316_IO_out, c0_n317_IO_out, c0_n318_IO_out, c0_n319_IO_out, c0_n320_IO_out, c0_n321_IO_out, c0_n322_IO_out, c0_n323_IO_out, c0_n324_IO_out, c0_n325_IO_out, c0_n326_IO_out, c0_n327_IO_out, c0_n328_IO_out, c0_n329_IO_out, c0_n330_IO_out, c0_n331_IO_out, c0_n332_IO_out, c0_n333_IO_out, c0_n334_IO_out, c0_n335_IO_out, c0_n336_IO_out, c0_n337_IO_out, c0_n338_IO_out, c0_n339_IO_out, c0_n340_IO_out, c0_n341_IO_out, c0_n342_IO_out, c0_n343_IO_out, c0_n344_IO_out, c0_n345_IO_out, c0_n346_IO_out, c0_n347_IO_out, c0_n348_IO_out, c0_n349_IO_out, c0_n350_IO_out, c0_n351_IO_out, c0_n352_IO_out, c0_n353_IO_out, c0_n354_IO_out, c0_n355_IO_out, c0_n356_IO_out, c0_n357_IO_out, c0_n358_IO_out, c0_n359_IO_out, c0_n360_IO_out, c0_n361_IO_out, c0_n362_IO_out, c0_n363_IO_out, c0_n364_IO_out, c0_n365_IO_out, c0_n366_IO_out, c0_n367_IO_out, c0_n368_IO_out, c0_n369_IO_out, c0_n370_IO_out, c0_n371_IO_out, c0_n372_IO_out, c0_n373_IO_out, c0_n374_IO_out, c0_n375_IO_out, c0_n376_IO_out, c0_n377_IO_out, c0_n378_IO_out, c0_n379_IO_out, c0_n380_IO_out, c0_n381_IO_out, c0_n382_IO_out, c0_n383_IO_out, c0_n384_IO_out, c0_n385_IO_out, c0_n386_IO_out, c0_n387_IO_out, c0_n388_IO_out, c0_n389_IO_out, c0_n390_IO_out, c0_n391_IO_out, c0_n392_IO_out, c0_n393_IO_out, c0_n394_IO_out, c0_n395_IO_out, c0_n396_IO_out, c0_n397_IO_out, c0_n398_IO_out, c0_n399_IO_out, c0_n400_IO_out, c0_n401_IO_out, c0_n402_IO_out, c0_n403_IO_out, c0_n404_IO_out, c0_n405_IO_out, c0_n406_IO_out, c0_n407_IO_out, c0_n408_IO_out, c0_n409_IO_out, c0_n410_IO_out, c0_n411_IO_out, c0_n412_IO_out, c0_n413_IO_out, c0_n414_IO_out, c0_n415_IO_out, c0_n416_IO_out, c0_n417_IO_out, c0_n418_IO_out, c0_n419_IO_out, c0_n420_IO_out, c0_n421_IO_out, c0_n422_IO_out, c0_n423_IO_out, c0_n424_IO_out, c0_n425_IO_out, c0_n426_IO_out, c0_n427_IO_out, c0_n428_IO_out, c0_n429_IO_out, c0_n430_IO_out, c0_n431_IO_out, c0_n432_IO_out, c0_n433_IO_out, c0_n434_IO_out, c0_n435_IO_out, c0_n436_IO_out, c0_n437_IO_out, c0_n438_IO_out, c0_n439_IO_out, c0_n440_IO_out, c0_n441_IO_out, c0_n442_IO_out, c0_n443_IO_out, c0_n444_IO_out, c0_n445_IO_out, c0_n446_IO_out, c0_n447_IO_out, c0_n448_IO_out, c0_n449_IO_out, c0_n450_IO_out, c0_n451_IO_out, c0_n452_IO_out, c0_n453_IO_out, c0_n454_IO_out, c0_n455_IO_out, c0_n456_IO_out, c0_n457_IO_out, c0_n458_IO_out, c0_n459_IO_out, c0_n460_IO_out, c0_n461_IO_out, c0_n462_IO_out, c0_n463_IO_out, c0_n464_IO_out, c0_n465_IO_out, c0_n466_IO_out, c0_n467_IO_out, c0_n468_IO_out, c0_n469_IO_out, c0_n470_IO_out, c0_n471_IO_out, c0_n472_IO_out, c0_n473_IO_out, c0_n474_IO_out, c0_n475_IO_out, c0_n476_IO_out, c0_n477_IO_out, c0_n478_IO_out, c0_n479_IO_out, c0_n480_IO_out, c0_n481_IO_out, c0_n482_IO_out, c0_n483_IO_out, c0_n484_IO_out, c0_n485_IO_out, c0_n486_IO_out, c0_n487_IO_out, c0_n488_IO_out, c0_n489_IO_out, c0_n490_IO_out, c0_n491_IO_out, c0_n492_IO_out, c0_n493_IO_out, c0_n494_IO_out, c0_n495_IO_out, c0_n496_IO_out, c0_n497_IO_out, c0_n498_IO_out, c0_n499_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c1_n0_IO_out, c1_n1_IO_out, c1_n2_IO_out, c1_n3_IO_out, c1_n4_IO_out, c1_n5_IO_out, c1_n6_IO_out, c1_n7_IO_out, c1_n8_IO_out, c1_n9_IO_out, c1_n10_IO_out, c1_n11_IO_out, c1_n12_IO_out, c1_n13_IO_out, c1_n14_IO_out, c1_n15_IO_out, c1_n16_IO_out, c1_n17_IO_out, c1_n18_IO_out, c1_n19_IO_out, c1_n20_IO_out, c1_n21_IO_out, c1_n22_IO_out, c1_n23_IO_out, c1_n24_IO_out, c1_n25_IO_out, c1_n26_IO_out, c1_n27_IO_out, c1_n28_IO_out, c1_n29_IO_out, c1_n30_IO_out, c1_n31_IO_out, c1_n32_IO_out, c1_n33_IO_out, c1_n34_IO_out, c1_n35_IO_out, c1_n36_IO_out, c1_n37_IO_out, c1_n38_IO_out, c1_n39_IO_out, c1_n40_IO_out, c1_n41_IO_out, c1_n42_IO_out, c1_n43_IO_out, c1_n44_IO_out, c1_n45_IO_out, c1_n46_IO_out, c1_n47_IO_out, c1_n48_IO_out, c1_n49_IO_out, c1_n50_IO_out, c1_n51_IO_out, c1_n52_IO_out, c1_n53_IO_out, c1_n54_IO_out, c1_n55_IO_out, c1_n56_IO_out, c1_n57_IO_out, c1_n58_IO_out, c1_n59_IO_out, c1_n60_IO_out, c1_n61_IO_out, c1_n62_IO_out, c1_n63_IO_out, c1_n64_IO_out, c1_n65_IO_out, c1_n66_IO_out, c1_n67_IO_out, c1_n68_IO_out, c1_n69_IO_out, c1_n70_IO_out, c1_n71_IO_out, c1_n72_IO_out, c1_n73_IO_out, c1_n74_IO_out, c1_n75_IO_out, c1_n76_IO_out, c1_n77_IO_out, c1_n78_IO_out, c1_n79_IO_out, c1_n80_IO_out, c1_n81_IO_out, c1_n82_IO_out, c1_n83_IO_out, c1_n84_IO_out, c1_n85_IO_out, c1_n86_IO_out, c1_n87_IO_out, c1_n88_IO_out, c1_n89_IO_out, c1_n90_IO_out, c1_n91_IO_out, c1_n92_IO_out, c1_n93_IO_out, c1_n94_IO_out, c1_n95_IO_out, c1_n96_IO_out, c1_n97_IO_out, c1_n98_IO_out, c1_n99_IO_out, c1_n100_IO_out, c1_n101_IO_out, c1_n102_IO_out, c1_n103_IO_out, c1_n104_IO_out, c1_n105_IO_out, c1_n106_IO_out, c1_n107_IO_out, c1_n108_IO_out, c1_n109_IO_out, c1_n110_IO_out, c1_n111_IO_out, c1_n112_IO_out, c1_n113_IO_out, c1_n114_IO_out, c1_n115_IO_out, c1_n116_IO_out, c1_n117_IO_out, c1_n118_IO_out, c1_n119_IO_out, c1_n120_IO_out, c1_n121_IO_out, c1_n122_IO_out, c1_n123_IO_out, c1_n124_IO_out, c1_n125_IO_out, c1_n126_IO_out, c1_n127_IO_out, c1_n128_IO_out, c1_n129_IO_out, c1_n130_IO_out, c1_n131_IO_out, c1_n132_IO_out, c1_n133_IO_out, c1_n134_IO_out, c1_n135_IO_out, c1_n136_IO_out, c1_n137_IO_out, c1_n138_IO_out, c1_n139_IO_out, c1_n140_IO_out, c1_n141_IO_out, c1_n142_IO_out, c1_n143_IO_out, c1_n144_IO_out, c1_n145_IO_out, c1_n146_IO_out, c1_n147_IO_out, c1_n148_IO_out, c1_n149_IO_out, c1_n150_IO_out, c1_n151_IO_out, c1_n152_IO_out, c1_n153_IO_out, c1_n154_IO_out, c1_n155_IO_out, c1_n156_IO_out, c1_n157_IO_out, c1_n158_IO_out, c1_n159_IO_out, c1_n160_IO_out, c1_n161_IO_out, c1_n162_IO_out, c1_n163_IO_out, c1_n164_IO_out, c1_n165_IO_out, c1_n166_IO_out, c1_n167_IO_out, c1_n168_IO_out, c1_n169_IO_out, c1_n170_IO_out, c1_n171_IO_out, c1_n172_IO_out, c1_n173_IO_out, c1_n174_IO_out, c1_n175_IO_out, c1_n176_IO_out, c1_n177_IO_out, c1_n178_IO_out, c1_n179_IO_out, c1_n180_IO_out, c1_n181_IO_out, c1_n182_IO_out, c1_n183_IO_out, c1_n184_IO_out, c1_n185_IO_out, c1_n186_IO_out, c1_n187_IO_out, c1_n188_IO_out, c1_n189_IO_out, c1_n190_IO_out, c1_n191_IO_out, c1_n192_IO_out, c1_n193_IO_out, c1_n194_IO_out, c1_n195_IO_out, c1_n196_IO_out, c1_n197_IO_out, c1_n198_IO_out, c1_n199_IO_out, c1_n200_IO_out, c1_n201_IO_out, c1_n202_IO_out, c1_n203_IO_out, c1_n204_IO_out, c1_n205_IO_out, c1_n206_IO_out, c1_n207_IO_out, c1_n208_IO_out, c1_n209_IO_out, c1_n210_IO_out, c1_n211_IO_out, c1_n212_IO_out, c1_n213_IO_out, c1_n214_IO_out, c1_n215_IO_out, c1_n216_IO_out, c1_n217_IO_out, c1_n218_IO_out, c1_n219_IO_out, c1_n220_IO_out, c1_n221_IO_out, c1_n222_IO_out, c1_n223_IO_out, c1_n224_IO_out, c1_n225_IO_out, c1_n226_IO_out, c1_n227_IO_out, c1_n228_IO_out, c1_n229_IO_out, c1_n230_IO_out, c1_n231_IO_out, c1_n232_IO_out, c1_n233_IO_out, c1_n234_IO_out, c1_n235_IO_out, c1_n236_IO_out, c1_n237_IO_out, c1_n238_IO_out, c1_n239_IO_out, c1_n240_IO_out, c1_n241_IO_out, c1_n242_IO_out, c1_n243_IO_out, c1_n244_IO_out, c1_n245_IO_out, c1_n246_IO_out, c1_n247_IO_out, c1_n248_IO_out, c1_n249_IO_out, c1_n250_IO_out, c1_n251_IO_out, c1_n252_IO_out, c1_n253_IO_out, c1_n254_IO_out, c1_n255_IO_out, c1_n256_IO_out, c1_n257_IO_out, c1_n258_IO_out, c1_n259_IO_out, c1_n260_IO_out, c1_n261_IO_out, c1_n262_IO_out, c1_n263_IO_out, c1_n264_IO_out, c1_n265_IO_out, c1_n266_IO_out, c1_n267_IO_out, c1_n268_IO_out, c1_n269_IO_out, c1_n270_IO_out, c1_n271_IO_out, c1_n272_IO_out, c1_n273_IO_out, c1_n274_IO_out, c1_n275_IO_out, c1_n276_IO_out, c1_n277_IO_out, c1_n278_IO_out, c1_n279_IO_out, c1_n280_IO_out, c1_n281_IO_out, c1_n282_IO_out, c1_n283_IO_out, c1_n284_IO_out, c1_n285_IO_out, c1_n286_IO_out, c1_n287_IO_out, c1_n288_IO_out, c1_n289_IO_out, c1_n290_IO_out, c1_n291_IO_out, c1_n292_IO_out, c1_n293_IO_out, c1_n294_IO_out, c1_n295_IO_out, c1_n296_IO_out, c1_n297_IO_out, c1_n298_IO_out, c1_n299_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c2_n0_IO_out, c2_n1_IO_out, c2_n2_IO_out, c2_n3_IO_out, c2_n4_IO_out, c2_n5_IO_out, c2_n6_IO_out, c2_n7_IO_out, c2_n8_IO_out, c2_n9_IO_out, c2_n10_IO_out, c2_n11_IO_out, c2_n12_IO_out, c2_n13_IO_out, c2_n14_IO_out, c2_n15_IO_out, c2_n16_IO_out, c2_n17_IO_out, c2_n18_IO_out, c2_n19_IO_out, c2_n20_IO_out, c2_n21_IO_out, c2_n22_IO_out, c2_n23_IO_out, c2_n24_IO_out, c2_n25_IO_out, c2_n26_IO_out, c2_n27_IO_out, c2_n28_IO_out, c2_n29_IO_out, c2_n30_IO_out, c2_n31_IO_out, c2_n32_IO_out, c2_n33_IO_out, c2_n34_IO_out, c2_n35_IO_out, c2_n36_IO_out, c2_n37_IO_out, c2_n38_IO_out, c2_n39_IO_out, c2_n40_IO_out, c2_n41_IO_out, c2_n42_IO_out, c2_n43_IO_out, c2_n44_IO_out, c2_n45_IO_out, c2_n46_IO_out, c2_n47_IO_out, c2_n48_IO_out, c2_n49_IO_out, c2_n50_IO_out, c2_n51_IO_out, c2_n52_IO_out, c2_n53_IO_out, c2_n54_IO_out, c2_n55_IO_out, c2_n56_IO_out, c2_n57_IO_out, c2_n58_IO_out, c2_n59_IO_out, c2_n60_IO_out, c2_n61_IO_out, c2_n62_IO_out, c2_n63_IO_out, c2_n64_IO_out, c2_n65_IO_out, c2_n66_IO_out, c2_n67_IO_out, c2_n68_IO_out, c2_n69_IO_out, c2_n70_IO_out, c2_n71_IO_out, c2_n72_IO_out, c2_n73_IO_out, c2_n74_IO_out, c2_n75_IO_out, c2_n76_IO_out, c2_n77_IO_out, c2_n78_IO_out, c2_n79_IO_out, c2_n80_IO_out, c2_n81_IO_out, c2_n82_IO_out, c2_n83_IO_out, c2_n84_IO_out, c2_n85_IO_out, c2_n86_IO_out, c2_n87_IO_out, c2_n88_IO_out, c2_n89_IO_out, c2_n90_IO_out, c2_n91_IO_out, c2_n92_IO_out, c2_n93_IO_out, c2_n94_IO_out, c2_n95_IO_out, c2_n96_IO_out, c2_n97_IO_out, c2_n98_IO_out, c2_n99_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c3_n0_IO_out, c3_n1_IO_out, c3_n2_IO_out, c3_n3_IO_out, c3_n4_IO_out, c3_n5_IO_out, c3_n6_IO_out, c3_n7_IO_out, c3_n8_IO_out, c3_n9_IO_out, c3_n10_IO_out, c3_n11_IO_out, c3_n12_IO_out, c3_n13_IO_out, c3_n14_IO_out, c3_n15_IO_out, c3_n16_IO_out, c3_n17_IO_out, c3_n18_IO_out, c3_n19_IO_out, c3_n20_IO_out, c3_n21_IO_out, c3_n22_IO_out, c3_n23_IO_out, c3_n24_IO_out, c3_n25_IO_out, c3_n26_IO_out, c3_n27_IO_out, c3_n28_IO_out, c3_n29_IO_out, c3_n30_IO_out, c3_n31_IO_out, c3_n32_IO_out, c3_n33_IO_out, c3_n34_IO_out, c3_n35_IO_out, c3_n36_IO_out, c3_n37_IO_out, c3_n38_IO_out, c3_n39_IO_out, c3_n40_IO_out, c3_n41_IO_out, c3_n42_IO_out, c3_n43_IO_out, c3_n44_IO_out, c3_n45_IO_out, c3_n46_IO_out, c3_n47_IO_out, c3_n48_IO_out, c3_n49_IO_out, c3_n50_IO_out, c3_n51_IO_out, c3_n52_IO_out, c3_n53_IO_out, c3_n54_IO_out, c3_n55_IO_out, c3_n56_IO_out, c3_n57_IO_out, c3_n58_IO_out, c3_n59_IO_out, c3_n60_IO_out, c3_n61_IO_out, c3_n62_IO_out, c3_n63_IO_out, c3_n64_IO_out, c3_n65_IO_out, c3_n66_IO_out, c3_n67_IO_out, c3_n68_IO_out, c3_n69_IO_out, c3_n70_IO_out, c3_n71_IO_out, c3_n72_IO_out, c3_n73_IO_out, c3_n74_IO_out, c3_n75_IO_out, c3_n76_IO_out, c3_n77_IO_out, c3_n78_IO_out, c3_n79_IO_out, c3_n80_IO_out, c3_n81_IO_out, c3_n82_IO_out, c3_n83_IO_out, c3_n84_IO_out, c3_n85_IO_out, c3_n86_IO_out, c3_n87_IO_out, c3_n88_IO_out, c3_n89_IO_out, c3_n90_IO_out, c3_n91_IO_out, c3_n92_IO_out, c3_n93_IO_out, c3_n94_IO_out, c3_n95_IO_out, c3_n96_IO_out, c3_n97_IO_out, c3_n98_IO_out, c3_n99_IO_out, c3_n100_IO_out, c3_n101_IO_out, c3_n102_IO_out, c3_n103_IO_out, c3_n104_IO_out, c3_n105_IO_out, c3_n106_IO_out, c3_n107_IO_out, c3_n108_IO_out, c3_n109_IO_out, c3_n110_IO_out, c3_n111_IO_out, c3_n112_IO_out, c3_n113_IO_out, c3_n114_IO_out, c3_n115_IO_out, c3_n116_IO_out, c3_n117_IO_out, c3_n118_IO_out, c3_n119_IO_out, c3_n120_IO_out, c3_n121_IO_out, c3_n122_IO_out, c3_n123_IO_out, c3_n124_IO_out, c3_n125_IO_out, c3_n126_IO_out, c3_n127_IO_out, c3_n128_IO_out, c3_n129_IO_out, c3_n130_IO_out, c3_n131_IO_out, c3_n132_IO_out, c3_n133_IO_out, c3_n134_IO_out, c3_n135_IO_out, c3_n136_IO_out, c3_n137_IO_out, c3_n138_IO_out, c3_n139_IO_out, c3_n140_IO_out, c3_n141_IO_out, c3_n142_IO_out, c3_n143_IO_out, c3_n144_IO_out, c3_n145_IO_out, c3_n146_IO_out, c3_n147_IO_out, c3_n148_IO_out, c3_n149_IO_out, c3_n150_IO_out, c3_n151_IO_out, c3_n152_IO_out, c3_n153_IO_out, c3_n154_IO_out, c3_n155_IO_out, c3_n156_IO_out, c3_n157_IO_out, c3_n158_IO_out, c3_n159_IO_out, c3_n160_IO_out, c3_n161_IO_out, c3_n162_IO_out, c3_n163_IO_out, c3_n164_IO_out, c3_n165_IO_out, c3_n166_IO_out, c3_n167_IO_out, c3_n168_IO_out, c3_n169_IO_out, c3_n170_IO_out, c3_n171_IO_out, c3_n172_IO_out, c3_n173_IO_out, c3_n174_IO_out, c3_n175_IO_out, c3_n176_IO_out, c3_n177_IO_out, c3_n178_IO_out, c3_n179_IO_out, c3_n180_IO_out, c3_n181_IO_out, c3_n182_IO_out, c3_n183_IO_out, c3_n184_IO_out, c3_n185_IO_out, c3_n186_IO_out, c3_n187_IO_out, c3_n188_IO_out, c3_n189_IO_out, c3_n190_IO_out, c3_n191_IO_out, c3_n192_IO_out, c3_n193_IO_out, c3_n194_IO_out, c3_n195_IO_out, c3_n196_IO_out, c3_n197_IO_out, c3_n198_IO_out, c3_n199_IO_out, c3_n200_IO_out, c3_n201_IO_out, c3_n202_IO_out, c3_n203_IO_out, c3_n204_IO_out, c3_n205_IO_out, c3_n206_IO_out, c3_n207_IO_out, c3_n208_IO_out, c3_n209_IO_out, c3_n210_IO_out, c3_n211_IO_out, c3_n212_IO_out, c3_n213_IO_out, c3_n214_IO_out, c3_n215_IO_out, c3_n216_IO_out, c3_n217_IO_out, c3_n218_IO_out, c3_n219_IO_out, c3_n220_IO_out, c3_n221_IO_out, c3_n222_IO_out, c3_n223_IO_out, c3_n224_IO_out, c3_n225_IO_out, c3_n226_IO_out, c3_n227_IO_out, c3_n228_IO_out, c3_n229_IO_out, c3_n230_IO_out, c3_n231_IO_out, c3_n232_IO_out, c3_n233_IO_out, c3_n234_IO_out, c3_n235_IO_out, c3_n236_IO_out, c3_n237_IO_out, c3_n238_IO_out, c3_n239_IO_out, c3_n240_IO_out, c3_n241_IO_out, c3_n242_IO_out, c3_n243_IO_out, c3_n244_IO_out, c3_n245_IO_out, c3_n246_IO_out, c3_n247_IO_out, c3_n248_IO_out, c3_n249_IO_out, c3_n250_IO_out, c3_n251_IO_out, c3_n252_IO_out, c3_n253_IO_out, c3_n254_IO_out, c3_n255_IO_out, c3_n256_IO_out, c3_n257_IO_out, c3_n258_IO_out, c3_n259_IO_out, c3_n260_IO_out, c3_n261_IO_out, c3_n262_IO_out, c3_n263_IO_out, c3_n264_IO_out, c3_n265_IO_out, c3_n266_IO_out, c3_n267_IO_out, c3_n268_IO_out, c3_n269_IO_out, c3_n270_IO_out, c3_n271_IO_out, c3_n272_IO_out, c3_n273_IO_out, c3_n274_IO_out, c3_n275_IO_out, c3_n276_IO_out, c3_n277_IO_out, c3_n278_IO_out, c3_n279_IO_out, c3_n280_IO_out, c3_n281_IO_out, c3_n282_IO_out, c3_n283_IO_out, c3_n284_IO_out, c3_n285_IO_out, c3_n286_IO_out, c3_n287_IO_out, c3_n288_IO_out, c3_n289_IO_out, c3_n290_IO_out, c3_n291_IO_out, c3_n292_IO_out, c3_n293_IO_out, c3_n294_IO_out, c3_n295_IO_out, c3_n296_IO_out, c3_n297_IO_out, c3_n298_IO_out, c3_n299_IO_out: SIGNED(BITS -1 DOWNTO 0);
    SIGNAL reg_IO_in: signed(TOTAL_BITS - 1 DOWNTO 0);
    SIGNAL en_registers: STD_LOGIC;
BEGIN
  en_registers <= update_weights AND clk;
  c1_IO_in <= c0_n0_IO_out & c0_n1_IO_out & c0_n2_IO_out & c0_n3_IO_out & c0_n4_IO_out & c0_n5_IO_out & c0_n6_IO_out & c0_n7_IO_out & c0_n8_IO_out & c0_n9_IO_out & c0_n10_IO_out & c0_n11_IO_out & c0_n12_IO_out & c0_n13_IO_out & c0_n14_IO_out & c0_n15_IO_out & c0_n16_IO_out & c0_n17_IO_out & c0_n18_IO_out & c0_n19_IO_out & c0_n20_IO_out & c0_n21_IO_out & c0_n22_IO_out & c0_n23_IO_out & c0_n24_IO_out & c0_n25_IO_out & c0_n26_IO_out & c0_n27_IO_out & c0_n28_IO_out & c0_n29_IO_out & c0_n30_IO_out & c0_n31_IO_out & c0_n32_IO_out & c0_n33_IO_out & c0_n34_IO_out & c0_n35_IO_out & c0_n36_IO_out & c0_n37_IO_out & c0_n38_IO_out & c0_n39_IO_out & c0_n40_IO_out & c0_n41_IO_out & c0_n42_IO_out & c0_n43_IO_out & c0_n44_IO_out & c0_n45_IO_out & c0_n46_IO_out & c0_n47_IO_out & c0_n48_IO_out & c0_n49_IO_out & c0_n50_IO_out & c0_n51_IO_out & c0_n52_IO_out & c0_n53_IO_out & c0_n54_IO_out & c0_n55_IO_out & c0_n56_IO_out & c0_n57_IO_out & c0_n58_IO_out & c0_n59_IO_out & c0_n60_IO_out & c0_n61_IO_out & c0_n62_IO_out & c0_n63_IO_out & c0_n64_IO_out & c0_n65_IO_out & c0_n66_IO_out & c0_n67_IO_out & c0_n68_IO_out & c0_n69_IO_out & c0_n70_IO_out & c0_n71_IO_out & c0_n72_IO_out & c0_n73_IO_out & c0_n74_IO_out & c0_n75_IO_out & c0_n76_IO_out & c0_n77_IO_out & c0_n78_IO_out & c0_n79_IO_out & c0_n80_IO_out & c0_n81_IO_out & c0_n82_IO_out & c0_n83_IO_out & c0_n84_IO_out & c0_n85_IO_out & c0_n86_IO_out & c0_n87_IO_out & c0_n88_IO_out & c0_n89_IO_out & c0_n90_IO_out & c0_n91_IO_out & c0_n92_IO_out & c0_n93_IO_out & c0_n94_IO_out & c0_n95_IO_out & c0_n96_IO_out & c0_n97_IO_out & c0_n98_IO_out & c0_n99_IO_out & c0_n100_IO_out & c0_n101_IO_out & c0_n102_IO_out & c0_n103_IO_out & c0_n104_IO_out & c0_n105_IO_out & c0_n106_IO_out & c0_n107_IO_out & c0_n108_IO_out & c0_n109_IO_out & c0_n110_IO_out & c0_n111_IO_out & c0_n112_IO_out & c0_n113_IO_out & c0_n114_IO_out & c0_n115_IO_out & c0_n116_IO_out & c0_n117_IO_out & c0_n118_IO_out & c0_n119_IO_out & c0_n120_IO_out & c0_n121_IO_out & c0_n122_IO_out & c0_n123_IO_out & c0_n124_IO_out & c0_n125_IO_out & c0_n126_IO_out & c0_n127_IO_out & c0_n128_IO_out & c0_n129_IO_out & c0_n130_IO_out & c0_n131_IO_out & c0_n132_IO_out & c0_n133_IO_out & c0_n134_IO_out & c0_n135_IO_out & c0_n136_IO_out & c0_n137_IO_out & c0_n138_IO_out & c0_n139_IO_out & c0_n140_IO_out & c0_n141_IO_out & c0_n142_IO_out & c0_n143_IO_out & c0_n144_IO_out & c0_n145_IO_out & c0_n146_IO_out & c0_n147_IO_out & c0_n148_IO_out & c0_n149_IO_out & c0_n150_IO_out & c0_n151_IO_out & c0_n152_IO_out & c0_n153_IO_out & c0_n154_IO_out & c0_n155_IO_out & c0_n156_IO_out & c0_n157_IO_out & c0_n158_IO_out & c0_n159_IO_out & c0_n160_IO_out & c0_n161_IO_out & c0_n162_IO_out & c0_n163_IO_out & c0_n164_IO_out & c0_n165_IO_out & c0_n166_IO_out & c0_n167_IO_out & c0_n168_IO_out & c0_n169_IO_out & c0_n170_IO_out & c0_n171_IO_out & c0_n172_IO_out & c0_n173_IO_out & c0_n174_IO_out & c0_n175_IO_out & c0_n176_IO_out & c0_n177_IO_out & c0_n178_IO_out & c0_n179_IO_out & c0_n180_IO_out & c0_n181_IO_out & c0_n182_IO_out & c0_n183_IO_out & c0_n184_IO_out & c0_n185_IO_out & c0_n186_IO_out & c0_n187_IO_out & c0_n188_IO_out & c0_n189_IO_out & c0_n190_IO_out & c0_n191_IO_out & c0_n192_IO_out & c0_n193_IO_out & c0_n194_IO_out & c0_n195_IO_out & c0_n196_IO_out & c0_n197_IO_out & c0_n198_IO_out & c0_n199_IO_out & c0_n200_IO_out & c0_n201_IO_out & c0_n202_IO_out & c0_n203_IO_out & c0_n204_IO_out & c0_n205_IO_out & c0_n206_IO_out & c0_n207_IO_out & c0_n208_IO_out & c0_n209_IO_out & c0_n210_IO_out & c0_n211_IO_out & c0_n212_IO_out & c0_n213_IO_out & c0_n214_IO_out & c0_n215_IO_out & c0_n216_IO_out & c0_n217_IO_out & c0_n218_IO_out & c0_n219_IO_out & c0_n220_IO_out & c0_n221_IO_out & c0_n222_IO_out & c0_n223_IO_out & c0_n224_IO_out & c0_n225_IO_out & c0_n226_IO_out & c0_n227_IO_out & c0_n228_IO_out & c0_n229_IO_out & c0_n230_IO_out & c0_n231_IO_out & c0_n232_IO_out & c0_n233_IO_out & c0_n234_IO_out & c0_n235_IO_out & c0_n236_IO_out & c0_n237_IO_out & c0_n238_IO_out & c0_n239_IO_out & c0_n240_IO_out & c0_n241_IO_out & c0_n242_IO_out & c0_n243_IO_out & c0_n244_IO_out & c0_n245_IO_out & c0_n246_IO_out & c0_n247_IO_out & c0_n248_IO_out & c0_n249_IO_out & c0_n250_IO_out & c0_n251_IO_out & c0_n252_IO_out & c0_n253_IO_out & c0_n254_IO_out & c0_n255_IO_out & c0_n256_IO_out & c0_n257_IO_out & c0_n258_IO_out & c0_n259_IO_out & c0_n260_IO_out & c0_n261_IO_out & c0_n262_IO_out & c0_n263_IO_out & c0_n264_IO_out & c0_n265_IO_out & c0_n266_IO_out & c0_n267_IO_out & c0_n268_IO_out & c0_n269_IO_out & c0_n270_IO_out & c0_n271_IO_out & c0_n272_IO_out & c0_n273_IO_out & c0_n274_IO_out & c0_n275_IO_out & c0_n276_IO_out & c0_n277_IO_out & c0_n278_IO_out & c0_n279_IO_out & c0_n280_IO_out & c0_n281_IO_out & c0_n282_IO_out & c0_n283_IO_out & c0_n284_IO_out & c0_n285_IO_out & c0_n286_IO_out & c0_n287_IO_out & c0_n288_IO_out & c0_n289_IO_out & c0_n290_IO_out & c0_n291_IO_out & c0_n292_IO_out & c0_n293_IO_out & c0_n294_IO_out & c0_n295_IO_out & c0_n296_IO_out & c0_n297_IO_out & c0_n298_IO_out & c0_n299_IO_out & c0_n300_IO_out & c0_n301_IO_out & c0_n302_IO_out & c0_n303_IO_out & c0_n304_IO_out & c0_n305_IO_out & c0_n306_IO_out & c0_n307_IO_out & c0_n308_IO_out & c0_n309_IO_out & c0_n310_IO_out & c0_n311_IO_out & c0_n312_IO_out & c0_n313_IO_out & c0_n314_IO_out & c0_n315_IO_out & c0_n316_IO_out & c0_n317_IO_out & c0_n318_IO_out & c0_n319_IO_out & c0_n320_IO_out & c0_n321_IO_out & c0_n322_IO_out & c0_n323_IO_out & c0_n324_IO_out & c0_n325_IO_out & c0_n326_IO_out & c0_n327_IO_out & c0_n328_IO_out & c0_n329_IO_out & c0_n330_IO_out & c0_n331_IO_out & c0_n332_IO_out & c0_n333_IO_out & c0_n334_IO_out & c0_n335_IO_out & c0_n336_IO_out & c0_n337_IO_out & c0_n338_IO_out & c0_n339_IO_out & c0_n340_IO_out & c0_n341_IO_out & c0_n342_IO_out & c0_n343_IO_out & c0_n344_IO_out & c0_n345_IO_out & c0_n346_IO_out & c0_n347_IO_out & c0_n348_IO_out & c0_n349_IO_out & c0_n350_IO_out & c0_n351_IO_out & c0_n352_IO_out & c0_n353_IO_out & c0_n354_IO_out & c0_n355_IO_out & c0_n356_IO_out & c0_n357_IO_out & c0_n358_IO_out & c0_n359_IO_out & c0_n360_IO_out & c0_n361_IO_out & c0_n362_IO_out & c0_n363_IO_out & c0_n364_IO_out & c0_n365_IO_out & c0_n366_IO_out & c0_n367_IO_out & c0_n368_IO_out & c0_n369_IO_out & c0_n370_IO_out & c0_n371_IO_out & c0_n372_IO_out & c0_n373_IO_out & c0_n374_IO_out & c0_n375_IO_out & c0_n376_IO_out & c0_n377_IO_out & c0_n378_IO_out & c0_n379_IO_out & c0_n380_IO_out & c0_n381_IO_out & c0_n382_IO_out & c0_n383_IO_out & c0_n384_IO_out & c0_n385_IO_out & c0_n386_IO_out & c0_n387_IO_out & c0_n388_IO_out & c0_n389_IO_out & c0_n390_IO_out & c0_n391_IO_out & c0_n392_IO_out & c0_n393_IO_out & c0_n394_IO_out & c0_n395_IO_out & c0_n396_IO_out & c0_n397_IO_out & c0_n398_IO_out & c0_n399_IO_out & c0_n400_IO_out & c0_n401_IO_out & c0_n402_IO_out & c0_n403_IO_out & c0_n404_IO_out & c0_n405_IO_out & c0_n406_IO_out & c0_n407_IO_out & c0_n408_IO_out & c0_n409_IO_out & c0_n410_IO_out & c0_n411_IO_out & c0_n412_IO_out & c0_n413_IO_out & c0_n414_IO_out & c0_n415_IO_out & c0_n416_IO_out & c0_n417_IO_out & c0_n418_IO_out & c0_n419_IO_out & c0_n420_IO_out & c0_n421_IO_out & c0_n422_IO_out & c0_n423_IO_out & c0_n424_IO_out & c0_n425_IO_out & c0_n426_IO_out & c0_n427_IO_out & c0_n428_IO_out & c0_n429_IO_out & c0_n430_IO_out & c0_n431_IO_out & c0_n432_IO_out & c0_n433_IO_out & c0_n434_IO_out & c0_n435_IO_out & c0_n436_IO_out & c0_n437_IO_out & c0_n438_IO_out & c0_n439_IO_out & c0_n440_IO_out & c0_n441_IO_out & c0_n442_IO_out & c0_n443_IO_out & c0_n444_IO_out & c0_n445_IO_out & c0_n446_IO_out & c0_n447_IO_out & c0_n448_IO_out & c0_n449_IO_out & c0_n450_IO_out & c0_n451_IO_out & c0_n452_IO_out & c0_n453_IO_out & c0_n454_IO_out & c0_n455_IO_out & c0_n456_IO_out & c0_n457_IO_out & c0_n458_IO_out & c0_n459_IO_out & c0_n460_IO_out & c0_n461_IO_out & c0_n462_IO_out & c0_n463_IO_out & c0_n464_IO_out & c0_n465_IO_out & c0_n466_IO_out & c0_n467_IO_out & c0_n468_IO_out & c0_n469_IO_out & c0_n470_IO_out & c0_n471_IO_out & c0_n472_IO_out & c0_n473_IO_out & c0_n474_IO_out & c0_n475_IO_out & c0_n476_IO_out & c0_n477_IO_out & c0_n478_IO_out & c0_n479_IO_out & c0_n480_IO_out & c0_n481_IO_out & c0_n482_IO_out & c0_n483_IO_out & c0_n484_IO_out & c0_n485_IO_out & c0_n486_IO_out & c0_n487_IO_out & c0_n488_IO_out & c0_n489_IO_out & c0_n490_IO_out & c0_n491_IO_out & c0_n492_IO_out & c0_n493_IO_out & c0_n494_IO_out & c0_n495_IO_out & c0_n496_IO_out & c0_n497_IO_out & c0_n498_IO_out & c0_n499_IO_out;
c2_IO_in <= c1_n0_IO_out & c1_n1_IO_out & c1_n2_IO_out & c1_n3_IO_out & c1_n4_IO_out & c1_n5_IO_out & c1_n6_IO_out & c1_n7_IO_out & c1_n8_IO_out & c1_n9_IO_out & c1_n10_IO_out & c1_n11_IO_out & c1_n12_IO_out & c1_n13_IO_out & c1_n14_IO_out & c1_n15_IO_out & c1_n16_IO_out & c1_n17_IO_out & c1_n18_IO_out & c1_n19_IO_out & c1_n20_IO_out & c1_n21_IO_out & c1_n22_IO_out & c1_n23_IO_out & c1_n24_IO_out & c1_n25_IO_out & c1_n26_IO_out & c1_n27_IO_out & c1_n28_IO_out & c1_n29_IO_out & c1_n30_IO_out & c1_n31_IO_out & c1_n32_IO_out & c1_n33_IO_out & c1_n34_IO_out & c1_n35_IO_out & c1_n36_IO_out & c1_n37_IO_out & c1_n38_IO_out & c1_n39_IO_out & c1_n40_IO_out & c1_n41_IO_out & c1_n42_IO_out & c1_n43_IO_out & c1_n44_IO_out & c1_n45_IO_out & c1_n46_IO_out & c1_n47_IO_out & c1_n48_IO_out & c1_n49_IO_out & c1_n50_IO_out & c1_n51_IO_out & c1_n52_IO_out & c1_n53_IO_out & c1_n54_IO_out & c1_n55_IO_out & c1_n56_IO_out & c1_n57_IO_out & c1_n58_IO_out & c1_n59_IO_out & c1_n60_IO_out & c1_n61_IO_out & c1_n62_IO_out & c1_n63_IO_out & c1_n64_IO_out & c1_n65_IO_out & c1_n66_IO_out & c1_n67_IO_out & c1_n68_IO_out & c1_n69_IO_out & c1_n70_IO_out & c1_n71_IO_out & c1_n72_IO_out & c1_n73_IO_out & c1_n74_IO_out & c1_n75_IO_out & c1_n76_IO_out & c1_n77_IO_out & c1_n78_IO_out & c1_n79_IO_out & c1_n80_IO_out & c1_n81_IO_out & c1_n82_IO_out & c1_n83_IO_out & c1_n84_IO_out & c1_n85_IO_out & c1_n86_IO_out & c1_n87_IO_out & c1_n88_IO_out & c1_n89_IO_out & c1_n90_IO_out & c1_n91_IO_out & c1_n92_IO_out & c1_n93_IO_out & c1_n94_IO_out & c1_n95_IO_out & c1_n96_IO_out & c1_n97_IO_out & c1_n98_IO_out & c1_n99_IO_out & c1_n100_IO_out & c1_n101_IO_out & c1_n102_IO_out & c1_n103_IO_out & c1_n104_IO_out & c1_n105_IO_out & c1_n106_IO_out & c1_n107_IO_out & c1_n108_IO_out & c1_n109_IO_out & c1_n110_IO_out & c1_n111_IO_out & c1_n112_IO_out & c1_n113_IO_out & c1_n114_IO_out & c1_n115_IO_out & c1_n116_IO_out & c1_n117_IO_out & c1_n118_IO_out & c1_n119_IO_out & c1_n120_IO_out & c1_n121_IO_out & c1_n122_IO_out & c1_n123_IO_out & c1_n124_IO_out & c1_n125_IO_out & c1_n126_IO_out & c1_n127_IO_out & c1_n128_IO_out & c1_n129_IO_out & c1_n130_IO_out & c1_n131_IO_out & c1_n132_IO_out & c1_n133_IO_out & c1_n134_IO_out & c1_n135_IO_out & c1_n136_IO_out & c1_n137_IO_out & c1_n138_IO_out & c1_n139_IO_out & c1_n140_IO_out & c1_n141_IO_out & c1_n142_IO_out & c1_n143_IO_out & c1_n144_IO_out & c1_n145_IO_out & c1_n146_IO_out & c1_n147_IO_out & c1_n148_IO_out & c1_n149_IO_out & c1_n150_IO_out & c1_n151_IO_out & c1_n152_IO_out & c1_n153_IO_out & c1_n154_IO_out & c1_n155_IO_out & c1_n156_IO_out & c1_n157_IO_out & c1_n158_IO_out & c1_n159_IO_out & c1_n160_IO_out & c1_n161_IO_out & c1_n162_IO_out & c1_n163_IO_out & c1_n164_IO_out & c1_n165_IO_out & c1_n166_IO_out & c1_n167_IO_out & c1_n168_IO_out & c1_n169_IO_out & c1_n170_IO_out & c1_n171_IO_out & c1_n172_IO_out & c1_n173_IO_out & c1_n174_IO_out & c1_n175_IO_out & c1_n176_IO_out & c1_n177_IO_out & c1_n178_IO_out & c1_n179_IO_out & c1_n180_IO_out & c1_n181_IO_out & c1_n182_IO_out & c1_n183_IO_out & c1_n184_IO_out & c1_n185_IO_out & c1_n186_IO_out & c1_n187_IO_out & c1_n188_IO_out & c1_n189_IO_out & c1_n190_IO_out & c1_n191_IO_out & c1_n192_IO_out & c1_n193_IO_out & c1_n194_IO_out & c1_n195_IO_out & c1_n196_IO_out & c1_n197_IO_out & c1_n198_IO_out & c1_n199_IO_out & c1_n200_IO_out & c1_n201_IO_out & c1_n202_IO_out & c1_n203_IO_out & c1_n204_IO_out & c1_n205_IO_out & c1_n206_IO_out & c1_n207_IO_out & c1_n208_IO_out & c1_n209_IO_out & c1_n210_IO_out & c1_n211_IO_out & c1_n212_IO_out & c1_n213_IO_out & c1_n214_IO_out & c1_n215_IO_out & c1_n216_IO_out & c1_n217_IO_out & c1_n218_IO_out & c1_n219_IO_out & c1_n220_IO_out & c1_n221_IO_out & c1_n222_IO_out & c1_n223_IO_out & c1_n224_IO_out & c1_n225_IO_out & c1_n226_IO_out & c1_n227_IO_out & c1_n228_IO_out & c1_n229_IO_out & c1_n230_IO_out & c1_n231_IO_out & c1_n232_IO_out & c1_n233_IO_out & c1_n234_IO_out & c1_n235_IO_out & c1_n236_IO_out & c1_n237_IO_out & c1_n238_IO_out & c1_n239_IO_out & c1_n240_IO_out & c1_n241_IO_out & c1_n242_IO_out & c1_n243_IO_out & c1_n244_IO_out & c1_n245_IO_out & c1_n246_IO_out & c1_n247_IO_out & c1_n248_IO_out & c1_n249_IO_out & c1_n250_IO_out & c1_n251_IO_out & c1_n252_IO_out & c1_n253_IO_out & c1_n254_IO_out & c1_n255_IO_out & c1_n256_IO_out & c1_n257_IO_out & c1_n258_IO_out & c1_n259_IO_out & c1_n260_IO_out & c1_n261_IO_out & c1_n262_IO_out & c1_n263_IO_out & c1_n264_IO_out & c1_n265_IO_out & c1_n266_IO_out & c1_n267_IO_out & c1_n268_IO_out & c1_n269_IO_out & c1_n270_IO_out & c1_n271_IO_out & c1_n272_IO_out & c1_n273_IO_out & c1_n274_IO_out & c1_n275_IO_out & c1_n276_IO_out & c1_n277_IO_out & c1_n278_IO_out & c1_n279_IO_out & c1_n280_IO_out & c1_n281_IO_out & c1_n282_IO_out & c1_n283_IO_out & c1_n284_IO_out & c1_n285_IO_out & c1_n286_IO_out & c1_n287_IO_out & c1_n288_IO_out & c1_n289_IO_out & c1_n290_IO_out & c1_n291_IO_out & c1_n292_IO_out & c1_n293_IO_out & c1_n294_IO_out & c1_n295_IO_out & c1_n296_IO_out & c1_n297_IO_out & c1_n298_IO_out & c1_n299_IO_out;
c3_IO_in <= c2_n0_IO_out & c2_n1_IO_out & c2_n2_IO_out & c2_n3_IO_out & c2_n4_IO_out & c2_n5_IO_out & c2_n6_IO_out & c2_n7_IO_out & c2_n8_IO_out & c2_n9_IO_out & c2_n10_IO_out & c2_n11_IO_out & c2_n12_IO_out & c2_n13_IO_out & c2_n14_IO_out & c2_n15_IO_out & c2_n16_IO_out & c2_n17_IO_out & c2_n18_IO_out & c2_n19_IO_out & c2_n20_IO_out & c2_n21_IO_out & c2_n22_IO_out & c2_n23_IO_out & c2_n24_IO_out & c2_n25_IO_out & c2_n26_IO_out & c2_n27_IO_out & c2_n28_IO_out & c2_n29_IO_out & c2_n30_IO_out & c2_n31_IO_out & c2_n32_IO_out & c2_n33_IO_out & c2_n34_IO_out & c2_n35_IO_out & c2_n36_IO_out & c2_n37_IO_out & c2_n38_IO_out & c2_n39_IO_out & c2_n40_IO_out & c2_n41_IO_out & c2_n42_IO_out & c2_n43_IO_out & c2_n44_IO_out & c2_n45_IO_out & c2_n46_IO_out & c2_n47_IO_out & c2_n48_IO_out & c2_n49_IO_out & c2_n50_IO_out & c2_n51_IO_out & c2_n52_IO_out & c2_n53_IO_out & c2_n54_IO_out & c2_n55_IO_out & c2_n56_IO_out & c2_n57_IO_out & c2_n58_IO_out & c2_n59_IO_out & c2_n60_IO_out & c2_n61_IO_out & c2_n62_IO_out & c2_n63_IO_out & c2_n64_IO_out & c2_n65_IO_out & c2_n66_IO_out & c2_n67_IO_out & c2_n68_IO_out & c2_n69_IO_out & c2_n70_IO_out & c2_n71_IO_out & c2_n72_IO_out & c2_n73_IO_out & c2_n74_IO_out & c2_n75_IO_out & c2_n76_IO_out & c2_n77_IO_out & c2_n78_IO_out & c2_n79_IO_out & c2_n80_IO_out & c2_n81_IO_out & c2_n82_IO_out & c2_n83_IO_out & c2_n84_IO_out & c2_n85_IO_out & c2_n86_IO_out & c2_n87_IO_out & c2_n88_IO_out & c2_n89_IO_out & c2_n90_IO_out & c2_n91_IO_out & c2_n92_IO_out & c2_n93_IO_out & c2_n94_IO_out & c2_n95_IO_out & c2_n96_IO_out & c2_n97_IO_out & c2_n98_IO_out & c2_n99_IO_out;
c4_IO_in <= c3_n0_IO_out & c3_n1_IO_out & c3_n2_IO_out & c3_n3_IO_out & c3_n4_IO_out & c3_n5_IO_out & c3_n6_IO_out & c3_n7_IO_out & c3_n8_IO_out & c3_n9_IO_out & c3_n10_IO_out & c3_n11_IO_out & c3_n12_IO_out & c3_n13_IO_out & c3_n14_IO_out & c3_n15_IO_out & c3_n16_IO_out & c3_n17_IO_out & c3_n18_IO_out & c3_n19_IO_out & c3_n20_IO_out & c3_n21_IO_out & c3_n22_IO_out & c3_n23_IO_out & c3_n24_IO_out & c3_n25_IO_out & c3_n26_IO_out & c3_n27_IO_out & c3_n28_IO_out & c3_n29_IO_out & c3_n30_IO_out & c3_n31_IO_out & c3_n32_IO_out & c3_n33_IO_out & c3_n34_IO_out & c3_n35_IO_out & c3_n36_IO_out & c3_n37_IO_out & c3_n38_IO_out & c3_n39_IO_out & c3_n40_IO_out & c3_n41_IO_out & c3_n42_IO_out & c3_n43_IO_out & c3_n44_IO_out & c3_n45_IO_out & c3_n46_IO_out & c3_n47_IO_out & c3_n48_IO_out & c3_n49_IO_out & c3_n50_IO_out & c3_n51_IO_out & c3_n52_IO_out & c3_n53_IO_out & c3_n54_IO_out & c3_n55_IO_out & c3_n56_IO_out & c3_n57_IO_out & c3_n58_IO_out & c3_n59_IO_out & c3_n60_IO_out & c3_n61_IO_out & c3_n62_IO_out & c3_n63_IO_out & c3_n64_IO_out & c3_n65_IO_out & c3_n66_IO_out & c3_n67_IO_out & c3_n68_IO_out & c3_n69_IO_out & c3_n70_IO_out & c3_n71_IO_out & c3_n72_IO_out & c3_n73_IO_out & c3_n74_IO_out & c3_n75_IO_out & c3_n76_IO_out & c3_n77_IO_out & c3_n78_IO_out & c3_n79_IO_out & c3_n80_IO_out & c3_n81_IO_out & c3_n82_IO_out & c3_n83_IO_out & c3_n84_IO_out & c3_n85_IO_out & c3_n86_IO_out & c3_n87_IO_out & c3_n88_IO_out & c3_n89_IO_out & c3_n90_IO_out & c3_n91_IO_out & c3_n92_IO_out & c3_n93_IO_out & c3_n94_IO_out & c3_n95_IO_out & c3_n96_IO_out & c3_n97_IO_out & c3_n98_IO_out & c3_n99_IO_out & c3_n100_IO_out & c3_n101_IO_out & c3_n102_IO_out & c3_n103_IO_out & c3_n104_IO_out & c3_n105_IO_out & c3_n106_IO_out & c3_n107_IO_out & c3_n108_IO_out & c3_n109_IO_out & c3_n110_IO_out & c3_n111_IO_out & c3_n112_IO_out & c3_n113_IO_out & c3_n114_IO_out & c3_n115_IO_out & c3_n116_IO_out & c3_n117_IO_out & c3_n118_IO_out & c3_n119_IO_out & c3_n120_IO_out & c3_n121_IO_out & c3_n122_IO_out & c3_n123_IO_out & c3_n124_IO_out & c3_n125_IO_out & c3_n126_IO_out & c3_n127_IO_out & c3_n128_IO_out & c3_n129_IO_out & c3_n130_IO_out & c3_n131_IO_out & c3_n132_IO_out & c3_n133_IO_out & c3_n134_IO_out & c3_n135_IO_out & c3_n136_IO_out & c3_n137_IO_out & c3_n138_IO_out & c3_n139_IO_out & c3_n140_IO_out & c3_n141_IO_out & c3_n142_IO_out & c3_n143_IO_out & c3_n144_IO_out & c3_n145_IO_out & c3_n146_IO_out & c3_n147_IO_out & c3_n148_IO_out & c3_n149_IO_out & c3_n150_IO_out & c3_n151_IO_out & c3_n152_IO_out & c3_n153_IO_out & c3_n154_IO_out & c3_n155_IO_out & c3_n156_IO_out & c3_n157_IO_out & c3_n158_IO_out & c3_n159_IO_out & c3_n160_IO_out & c3_n161_IO_out & c3_n162_IO_out & c3_n163_IO_out & c3_n164_IO_out & c3_n165_IO_out & c3_n166_IO_out & c3_n167_IO_out & c3_n168_IO_out & c3_n169_IO_out & c3_n170_IO_out & c3_n171_IO_out & c3_n172_IO_out & c3_n173_IO_out & c3_n174_IO_out & c3_n175_IO_out & c3_n176_IO_out & c3_n177_IO_out & c3_n178_IO_out & c3_n179_IO_out & c3_n180_IO_out & c3_n181_IO_out & c3_n182_IO_out & c3_n183_IO_out & c3_n184_IO_out & c3_n185_IO_out & c3_n186_IO_out & c3_n187_IO_out & c3_n188_IO_out & c3_n189_IO_out & c3_n190_IO_out & c3_n191_IO_out & c3_n192_IO_out & c3_n193_IO_out & c3_n194_IO_out & c3_n195_IO_out & c3_n196_IO_out & c3_n197_IO_out & c3_n198_IO_out & c3_n199_IO_out & c3_n200_IO_out & c3_n201_IO_out & c3_n202_IO_out & c3_n203_IO_out & c3_n204_IO_out & c3_n205_IO_out & c3_n206_IO_out & c3_n207_IO_out & c3_n208_IO_out & c3_n209_IO_out & c3_n210_IO_out & c3_n211_IO_out & c3_n212_IO_out & c3_n213_IO_out & c3_n214_IO_out & c3_n215_IO_out & c3_n216_IO_out & c3_n217_IO_out & c3_n218_IO_out & c3_n219_IO_out & c3_n220_IO_out & c3_n221_IO_out & c3_n222_IO_out & c3_n223_IO_out & c3_n224_IO_out & c3_n225_IO_out & c3_n226_IO_out & c3_n227_IO_out & c3_n228_IO_out & c3_n229_IO_out & c3_n230_IO_out & c3_n231_IO_out & c3_n232_IO_out & c3_n233_IO_out & c3_n234_IO_out & c3_n235_IO_out & c3_n236_IO_out & c3_n237_IO_out & c3_n238_IO_out & c3_n239_IO_out & c3_n240_IO_out & c3_n241_IO_out & c3_n242_IO_out & c3_n243_IO_out & c3_n244_IO_out & c3_n245_IO_out & c3_n246_IO_out & c3_n247_IO_out & c3_n248_IO_out & c3_n249_IO_out & c3_n250_IO_out & c3_n251_IO_out & c3_n252_IO_out & c3_n253_IO_out & c3_n254_IO_out & c3_n255_IO_out & c3_n256_IO_out & c3_n257_IO_out & c3_n258_IO_out & c3_n259_IO_out & c3_n260_IO_out & c3_n261_IO_out & c3_n262_IO_out & c3_n263_IO_out & c3_n264_IO_out & c3_n265_IO_out & c3_n266_IO_out & c3_n267_IO_out & c3_n268_IO_out & c3_n269_IO_out & c3_n270_IO_out & c3_n271_IO_out & c3_n272_IO_out & c3_n273_IO_out & c3_n274_IO_out & c3_n275_IO_out & c3_n276_IO_out & c3_n277_IO_out & c3_n278_IO_out & c3_n279_IO_out & c3_n280_IO_out & c3_n281_IO_out & c3_n282_IO_out & c3_n283_IO_out & c3_n284_IO_out & c3_n285_IO_out & c3_n286_IO_out & c3_n287_IO_out & c3_n288_IO_out & c3_n289_IO_out & c3_n290_IO_out & c3_n291_IO_out & c3_n292_IO_out & c3_n293_IO_out & c3_n294_IO_out & c3_n295_IO_out & c3_n296_IO_out & c3_n297_IO_out & c3_n298_IO_out & c3_n299_IO_out;

  PROCESS (clk, rst)
  BEGIN
    IF rst = '1' THEN
      reg_IO_in <= (OTHERS => '0');
    ELSIF clk'event AND clk = '1' THEN
      reg_IO_in <= IO_in;
    END IF;
  END PROCESS;

camada0_inst_0: ENTITY work.camada0_ReLU_500neuron_8bits_784n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> reg_IO_in, 
            c0_n0_W_in=> c0_n0_W_in, 
            c0_n1_W_in=> c0_n1_W_in, 
            c0_n2_W_in=> c0_n2_W_in, 
            c0_n3_W_in=> c0_n3_W_in, 
            c0_n4_W_in=> c0_n4_W_in, 
            c0_n5_W_in=> c0_n5_W_in, 
            c0_n6_W_in=> c0_n6_W_in, 
            c0_n7_W_in=> c0_n7_W_in, 
            c0_n8_W_in=> c0_n8_W_in, 
            c0_n9_W_in=> c0_n9_W_in, 
            c0_n10_W_in=> c0_n10_W_in, 
            c0_n11_W_in=> c0_n11_W_in, 
            c0_n12_W_in=> c0_n12_W_in, 
            c0_n13_W_in=> c0_n13_W_in, 
            c0_n14_W_in=> c0_n14_W_in, 
            c0_n15_W_in=> c0_n15_W_in, 
            c0_n16_W_in=> c0_n16_W_in, 
            c0_n17_W_in=> c0_n17_W_in, 
            c0_n18_W_in=> c0_n18_W_in, 
            c0_n19_W_in=> c0_n19_W_in, 
            c0_n20_W_in=> c0_n20_W_in, 
            c0_n21_W_in=> c0_n21_W_in, 
            c0_n22_W_in=> c0_n22_W_in, 
            c0_n23_W_in=> c0_n23_W_in, 
            c0_n24_W_in=> c0_n24_W_in, 
            c0_n25_W_in=> c0_n25_W_in, 
            c0_n26_W_in=> c0_n26_W_in, 
            c0_n27_W_in=> c0_n27_W_in, 
            c0_n28_W_in=> c0_n28_W_in, 
            c0_n29_W_in=> c0_n29_W_in, 
            c0_n30_W_in=> c0_n30_W_in, 
            c0_n31_W_in=> c0_n31_W_in, 
            c0_n32_W_in=> c0_n32_W_in, 
            c0_n33_W_in=> c0_n33_W_in, 
            c0_n34_W_in=> c0_n34_W_in, 
            c0_n35_W_in=> c0_n35_W_in, 
            c0_n36_W_in=> c0_n36_W_in, 
            c0_n37_W_in=> c0_n37_W_in, 
            c0_n38_W_in=> c0_n38_W_in, 
            c0_n39_W_in=> c0_n39_W_in, 
            c0_n40_W_in=> c0_n40_W_in, 
            c0_n41_W_in=> c0_n41_W_in, 
            c0_n42_W_in=> c0_n42_W_in, 
            c0_n43_W_in=> c0_n43_W_in, 
            c0_n44_W_in=> c0_n44_W_in, 
            c0_n45_W_in=> c0_n45_W_in, 
            c0_n46_W_in=> c0_n46_W_in, 
            c0_n47_W_in=> c0_n47_W_in, 
            c0_n48_W_in=> c0_n48_W_in, 
            c0_n49_W_in=> c0_n49_W_in, 
            c0_n50_W_in=> c0_n50_W_in, 
            c0_n51_W_in=> c0_n51_W_in, 
            c0_n52_W_in=> c0_n52_W_in, 
            c0_n53_W_in=> c0_n53_W_in, 
            c0_n54_W_in=> c0_n54_W_in, 
            c0_n55_W_in=> c0_n55_W_in, 
            c0_n56_W_in=> c0_n56_W_in, 
            c0_n57_W_in=> c0_n57_W_in, 
            c0_n58_W_in=> c0_n58_W_in, 
            c0_n59_W_in=> c0_n59_W_in, 
            c0_n60_W_in=> c0_n60_W_in, 
            c0_n61_W_in=> c0_n61_W_in, 
            c0_n62_W_in=> c0_n62_W_in, 
            c0_n63_W_in=> c0_n63_W_in, 
            c0_n64_W_in=> c0_n64_W_in, 
            c0_n65_W_in=> c0_n65_W_in, 
            c0_n66_W_in=> c0_n66_W_in, 
            c0_n67_W_in=> c0_n67_W_in, 
            c0_n68_W_in=> c0_n68_W_in, 
            c0_n69_W_in=> c0_n69_W_in, 
            c0_n70_W_in=> c0_n70_W_in, 
            c0_n71_W_in=> c0_n71_W_in, 
            c0_n72_W_in=> c0_n72_W_in, 
            c0_n73_W_in=> c0_n73_W_in, 
            c0_n74_W_in=> c0_n74_W_in, 
            c0_n75_W_in=> c0_n75_W_in, 
            c0_n76_W_in=> c0_n76_W_in, 
            c0_n77_W_in=> c0_n77_W_in, 
            c0_n78_W_in=> c0_n78_W_in, 
            c0_n79_W_in=> c0_n79_W_in, 
            c0_n80_W_in=> c0_n80_W_in, 
            c0_n81_W_in=> c0_n81_W_in, 
            c0_n82_W_in=> c0_n82_W_in, 
            c0_n83_W_in=> c0_n83_W_in, 
            c0_n84_W_in=> c0_n84_W_in, 
            c0_n85_W_in=> c0_n85_W_in, 
            c0_n86_W_in=> c0_n86_W_in, 
            c0_n87_W_in=> c0_n87_W_in, 
            c0_n88_W_in=> c0_n88_W_in, 
            c0_n89_W_in=> c0_n89_W_in, 
            c0_n90_W_in=> c0_n90_W_in, 
            c0_n91_W_in=> c0_n91_W_in, 
            c0_n92_W_in=> c0_n92_W_in, 
            c0_n93_W_in=> c0_n93_W_in, 
            c0_n94_W_in=> c0_n94_W_in, 
            c0_n95_W_in=> c0_n95_W_in, 
            c0_n96_W_in=> c0_n96_W_in, 
            c0_n97_W_in=> c0_n97_W_in, 
            c0_n98_W_in=> c0_n98_W_in, 
            c0_n99_W_in=> c0_n99_W_in, 
            c0_n100_W_in=> c0_n100_W_in, 
            c0_n101_W_in=> c0_n101_W_in, 
            c0_n102_W_in=> c0_n102_W_in, 
            c0_n103_W_in=> c0_n103_W_in, 
            c0_n104_W_in=> c0_n104_W_in, 
            c0_n105_W_in=> c0_n105_W_in, 
            c0_n106_W_in=> c0_n106_W_in, 
            c0_n107_W_in=> c0_n107_W_in, 
            c0_n108_W_in=> c0_n108_W_in, 
            c0_n109_W_in=> c0_n109_W_in, 
            c0_n110_W_in=> c0_n110_W_in, 
            c0_n111_W_in=> c0_n111_W_in, 
            c0_n112_W_in=> c0_n112_W_in, 
            c0_n113_W_in=> c0_n113_W_in, 
            c0_n114_W_in=> c0_n114_W_in, 
            c0_n115_W_in=> c0_n115_W_in, 
            c0_n116_W_in=> c0_n116_W_in, 
            c0_n117_W_in=> c0_n117_W_in, 
            c0_n118_W_in=> c0_n118_W_in, 
            c0_n119_W_in=> c0_n119_W_in, 
            c0_n120_W_in=> c0_n120_W_in, 
            c0_n121_W_in=> c0_n121_W_in, 
            c0_n122_W_in=> c0_n122_W_in, 
            c0_n123_W_in=> c0_n123_W_in, 
            c0_n124_W_in=> c0_n124_W_in, 
            c0_n125_W_in=> c0_n125_W_in, 
            c0_n126_W_in=> c0_n126_W_in, 
            c0_n127_W_in=> c0_n127_W_in, 
            c0_n128_W_in=> c0_n128_W_in, 
            c0_n129_W_in=> c0_n129_W_in, 
            c0_n130_W_in=> c0_n130_W_in, 
            c0_n131_W_in=> c0_n131_W_in, 
            c0_n132_W_in=> c0_n132_W_in, 
            c0_n133_W_in=> c0_n133_W_in, 
            c0_n134_W_in=> c0_n134_W_in, 
            c0_n135_W_in=> c0_n135_W_in, 
            c0_n136_W_in=> c0_n136_W_in, 
            c0_n137_W_in=> c0_n137_W_in, 
            c0_n138_W_in=> c0_n138_W_in, 
            c0_n139_W_in=> c0_n139_W_in, 
            c0_n140_W_in=> c0_n140_W_in, 
            c0_n141_W_in=> c0_n141_W_in, 
            c0_n142_W_in=> c0_n142_W_in, 
            c0_n143_W_in=> c0_n143_W_in, 
            c0_n144_W_in=> c0_n144_W_in, 
            c0_n145_W_in=> c0_n145_W_in, 
            c0_n146_W_in=> c0_n146_W_in, 
            c0_n147_W_in=> c0_n147_W_in, 
            c0_n148_W_in=> c0_n148_W_in, 
            c0_n149_W_in=> c0_n149_W_in, 
            c0_n150_W_in=> c0_n150_W_in, 
            c0_n151_W_in=> c0_n151_W_in, 
            c0_n152_W_in=> c0_n152_W_in, 
            c0_n153_W_in=> c0_n153_W_in, 
            c0_n154_W_in=> c0_n154_W_in, 
            c0_n155_W_in=> c0_n155_W_in, 
            c0_n156_W_in=> c0_n156_W_in, 
            c0_n157_W_in=> c0_n157_W_in, 
            c0_n158_W_in=> c0_n158_W_in, 
            c0_n159_W_in=> c0_n159_W_in, 
            c0_n160_W_in=> c0_n160_W_in, 
            c0_n161_W_in=> c0_n161_W_in, 
            c0_n162_W_in=> c0_n162_W_in, 
            c0_n163_W_in=> c0_n163_W_in, 
            c0_n164_W_in=> c0_n164_W_in, 
            c0_n165_W_in=> c0_n165_W_in, 
            c0_n166_W_in=> c0_n166_W_in, 
            c0_n167_W_in=> c0_n167_W_in, 
            c0_n168_W_in=> c0_n168_W_in, 
            c0_n169_W_in=> c0_n169_W_in, 
            c0_n170_W_in=> c0_n170_W_in, 
            c0_n171_W_in=> c0_n171_W_in, 
            c0_n172_W_in=> c0_n172_W_in, 
            c0_n173_W_in=> c0_n173_W_in, 
            c0_n174_W_in=> c0_n174_W_in, 
            c0_n175_W_in=> c0_n175_W_in, 
            c0_n176_W_in=> c0_n176_W_in, 
            c0_n177_W_in=> c0_n177_W_in, 
            c0_n178_W_in=> c0_n178_W_in, 
            c0_n179_W_in=> c0_n179_W_in, 
            c0_n180_W_in=> c0_n180_W_in, 
            c0_n181_W_in=> c0_n181_W_in, 
            c0_n182_W_in=> c0_n182_W_in, 
            c0_n183_W_in=> c0_n183_W_in, 
            c0_n184_W_in=> c0_n184_W_in, 
            c0_n185_W_in=> c0_n185_W_in, 
            c0_n186_W_in=> c0_n186_W_in, 
            c0_n187_W_in=> c0_n187_W_in, 
            c0_n188_W_in=> c0_n188_W_in, 
            c0_n189_W_in=> c0_n189_W_in, 
            c0_n190_W_in=> c0_n190_W_in, 
            c0_n191_W_in=> c0_n191_W_in, 
            c0_n192_W_in=> c0_n192_W_in, 
            c0_n193_W_in=> c0_n193_W_in, 
            c0_n194_W_in=> c0_n194_W_in, 
            c0_n195_W_in=> c0_n195_W_in, 
            c0_n196_W_in=> c0_n196_W_in, 
            c0_n197_W_in=> c0_n197_W_in, 
            c0_n198_W_in=> c0_n198_W_in, 
            c0_n199_W_in=> c0_n199_W_in, 
            c0_n200_W_in=> c0_n200_W_in, 
            c0_n201_W_in=> c0_n201_W_in, 
            c0_n202_W_in=> c0_n202_W_in, 
            c0_n203_W_in=> c0_n203_W_in, 
            c0_n204_W_in=> c0_n204_W_in, 
            c0_n205_W_in=> c0_n205_W_in, 
            c0_n206_W_in=> c0_n206_W_in, 
            c0_n207_W_in=> c0_n207_W_in, 
            c0_n208_W_in=> c0_n208_W_in, 
            c0_n209_W_in=> c0_n209_W_in, 
            c0_n210_W_in=> c0_n210_W_in, 
            c0_n211_W_in=> c0_n211_W_in, 
            c0_n212_W_in=> c0_n212_W_in, 
            c0_n213_W_in=> c0_n213_W_in, 
            c0_n214_W_in=> c0_n214_W_in, 
            c0_n215_W_in=> c0_n215_W_in, 
            c0_n216_W_in=> c0_n216_W_in, 
            c0_n217_W_in=> c0_n217_W_in, 
            c0_n218_W_in=> c0_n218_W_in, 
            c0_n219_W_in=> c0_n219_W_in, 
            c0_n220_W_in=> c0_n220_W_in, 
            c0_n221_W_in=> c0_n221_W_in, 
            c0_n222_W_in=> c0_n222_W_in, 
            c0_n223_W_in=> c0_n223_W_in, 
            c0_n224_W_in=> c0_n224_W_in, 
            c0_n225_W_in=> c0_n225_W_in, 
            c0_n226_W_in=> c0_n226_W_in, 
            c0_n227_W_in=> c0_n227_W_in, 
            c0_n228_W_in=> c0_n228_W_in, 
            c0_n229_W_in=> c0_n229_W_in, 
            c0_n230_W_in=> c0_n230_W_in, 
            c0_n231_W_in=> c0_n231_W_in, 
            c0_n232_W_in=> c0_n232_W_in, 
            c0_n233_W_in=> c0_n233_W_in, 
            c0_n234_W_in=> c0_n234_W_in, 
            c0_n235_W_in=> c0_n235_W_in, 
            c0_n236_W_in=> c0_n236_W_in, 
            c0_n237_W_in=> c0_n237_W_in, 
            c0_n238_W_in=> c0_n238_W_in, 
            c0_n239_W_in=> c0_n239_W_in, 
            c0_n240_W_in=> c0_n240_W_in, 
            c0_n241_W_in=> c0_n241_W_in, 
            c0_n242_W_in=> c0_n242_W_in, 
            c0_n243_W_in=> c0_n243_W_in, 
            c0_n244_W_in=> c0_n244_W_in, 
            c0_n245_W_in=> c0_n245_W_in, 
            c0_n246_W_in=> c0_n246_W_in, 
            c0_n247_W_in=> c0_n247_W_in, 
            c0_n248_W_in=> c0_n248_W_in, 
            c0_n249_W_in=> c0_n249_W_in, 
            c0_n250_W_in=> c0_n250_W_in, 
            c0_n251_W_in=> c0_n251_W_in, 
            c0_n252_W_in=> c0_n252_W_in, 
            c0_n253_W_in=> c0_n253_W_in, 
            c0_n254_W_in=> c0_n254_W_in, 
            c0_n255_W_in=> c0_n255_W_in, 
            c0_n256_W_in=> c0_n256_W_in, 
            c0_n257_W_in=> c0_n257_W_in, 
            c0_n258_W_in=> c0_n258_W_in, 
            c0_n259_W_in=> c0_n259_W_in, 
            c0_n260_W_in=> c0_n260_W_in, 
            c0_n261_W_in=> c0_n261_W_in, 
            c0_n262_W_in=> c0_n262_W_in, 
            c0_n263_W_in=> c0_n263_W_in, 
            c0_n264_W_in=> c0_n264_W_in, 
            c0_n265_W_in=> c0_n265_W_in, 
            c0_n266_W_in=> c0_n266_W_in, 
            c0_n267_W_in=> c0_n267_W_in, 
            c0_n268_W_in=> c0_n268_W_in, 
            c0_n269_W_in=> c0_n269_W_in, 
            c0_n270_W_in=> c0_n270_W_in, 
            c0_n271_W_in=> c0_n271_W_in, 
            c0_n272_W_in=> c0_n272_W_in, 
            c0_n273_W_in=> c0_n273_W_in, 
            c0_n274_W_in=> c0_n274_W_in, 
            c0_n275_W_in=> c0_n275_W_in, 
            c0_n276_W_in=> c0_n276_W_in, 
            c0_n277_W_in=> c0_n277_W_in, 
            c0_n278_W_in=> c0_n278_W_in, 
            c0_n279_W_in=> c0_n279_W_in, 
            c0_n280_W_in=> c0_n280_W_in, 
            c0_n281_W_in=> c0_n281_W_in, 
            c0_n282_W_in=> c0_n282_W_in, 
            c0_n283_W_in=> c0_n283_W_in, 
            c0_n284_W_in=> c0_n284_W_in, 
            c0_n285_W_in=> c0_n285_W_in, 
            c0_n286_W_in=> c0_n286_W_in, 
            c0_n287_W_in=> c0_n287_W_in, 
            c0_n288_W_in=> c0_n288_W_in, 
            c0_n289_W_in=> c0_n289_W_in, 
            c0_n290_W_in=> c0_n290_W_in, 
            c0_n291_W_in=> c0_n291_W_in, 
            c0_n292_W_in=> c0_n292_W_in, 
            c0_n293_W_in=> c0_n293_W_in, 
            c0_n294_W_in=> c0_n294_W_in, 
            c0_n295_W_in=> c0_n295_W_in, 
            c0_n296_W_in=> c0_n296_W_in, 
            c0_n297_W_in=> c0_n297_W_in, 
            c0_n298_W_in=> c0_n298_W_in, 
            c0_n299_W_in=> c0_n299_W_in, 
            c0_n300_W_in=> c0_n300_W_in, 
            c0_n301_W_in=> c0_n301_W_in, 
            c0_n302_W_in=> c0_n302_W_in, 
            c0_n303_W_in=> c0_n303_W_in, 
            c0_n304_W_in=> c0_n304_W_in, 
            c0_n305_W_in=> c0_n305_W_in, 
            c0_n306_W_in=> c0_n306_W_in, 
            c0_n307_W_in=> c0_n307_W_in, 
            c0_n308_W_in=> c0_n308_W_in, 
            c0_n309_W_in=> c0_n309_W_in, 
            c0_n310_W_in=> c0_n310_W_in, 
            c0_n311_W_in=> c0_n311_W_in, 
            c0_n312_W_in=> c0_n312_W_in, 
            c0_n313_W_in=> c0_n313_W_in, 
            c0_n314_W_in=> c0_n314_W_in, 
            c0_n315_W_in=> c0_n315_W_in, 
            c0_n316_W_in=> c0_n316_W_in, 
            c0_n317_W_in=> c0_n317_W_in, 
            c0_n318_W_in=> c0_n318_W_in, 
            c0_n319_W_in=> c0_n319_W_in, 
            c0_n320_W_in=> c0_n320_W_in, 
            c0_n321_W_in=> c0_n321_W_in, 
            c0_n322_W_in=> c0_n322_W_in, 
            c0_n323_W_in=> c0_n323_W_in, 
            c0_n324_W_in=> c0_n324_W_in, 
            c0_n325_W_in=> c0_n325_W_in, 
            c0_n326_W_in=> c0_n326_W_in, 
            c0_n327_W_in=> c0_n327_W_in, 
            c0_n328_W_in=> c0_n328_W_in, 
            c0_n329_W_in=> c0_n329_W_in, 
            c0_n330_W_in=> c0_n330_W_in, 
            c0_n331_W_in=> c0_n331_W_in, 
            c0_n332_W_in=> c0_n332_W_in, 
            c0_n333_W_in=> c0_n333_W_in, 
            c0_n334_W_in=> c0_n334_W_in, 
            c0_n335_W_in=> c0_n335_W_in, 
            c0_n336_W_in=> c0_n336_W_in, 
            c0_n337_W_in=> c0_n337_W_in, 
            c0_n338_W_in=> c0_n338_W_in, 
            c0_n339_W_in=> c0_n339_W_in, 
            c0_n340_W_in=> c0_n340_W_in, 
            c0_n341_W_in=> c0_n341_W_in, 
            c0_n342_W_in=> c0_n342_W_in, 
            c0_n343_W_in=> c0_n343_W_in, 
            c0_n344_W_in=> c0_n344_W_in, 
            c0_n345_W_in=> c0_n345_W_in, 
            c0_n346_W_in=> c0_n346_W_in, 
            c0_n347_W_in=> c0_n347_W_in, 
            c0_n348_W_in=> c0_n348_W_in, 
            c0_n349_W_in=> c0_n349_W_in, 
            c0_n350_W_in=> c0_n350_W_in, 
            c0_n351_W_in=> c0_n351_W_in, 
            c0_n352_W_in=> c0_n352_W_in, 
            c0_n353_W_in=> c0_n353_W_in, 
            c0_n354_W_in=> c0_n354_W_in, 
            c0_n355_W_in=> c0_n355_W_in, 
            c0_n356_W_in=> c0_n356_W_in, 
            c0_n357_W_in=> c0_n357_W_in, 
            c0_n358_W_in=> c0_n358_W_in, 
            c0_n359_W_in=> c0_n359_W_in, 
            c0_n360_W_in=> c0_n360_W_in, 
            c0_n361_W_in=> c0_n361_W_in, 
            c0_n362_W_in=> c0_n362_W_in, 
            c0_n363_W_in=> c0_n363_W_in, 
            c0_n364_W_in=> c0_n364_W_in, 
            c0_n365_W_in=> c0_n365_W_in, 
            c0_n366_W_in=> c0_n366_W_in, 
            c0_n367_W_in=> c0_n367_W_in, 
            c0_n368_W_in=> c0_n368_W_in, 
            c0_n369_W_in=> c0_n369_W_in, 
            c0_n370_W_in=> c0_n370_W_in, 
            c0_n371_W_in=> c0_n371_W_in, 
            c0_n372_W_in=> c0_n372_W_in, 
            c0_n373_W_in=> c0_n373_W_in, 
            c0_n374_W_in=> c0_n374_W_in, 
            c0_n375_W_in=> c0_n375_W_in, 
            c0_n376_W_in=> c0_n376_W_in, 
            c0_n377_W_in=> c0_n377_W_in, 
            c0_n378_W_in=> c0_n378_W_in, 
            c0_n379_W_in=> c0_n379_W_in, 
            c0_n380_W_in=> c0_n380_W_in, 
            c0_n381_W_in=> c0_n381_W_in, 
            c0_n382_W_in=> c0_n382_W_in, 
            c0_n383_W_in=> c0_n383_W_in, 
            c0_n384_W_in=> c0_n384_W_in, 
            c0_n385_W_in=> c0_n385_W_in, 
            c0_n386_W_in=> c0_n386_W_in, 
            c0_n387_W_in=> c0_n387_W_in, 
            c0_n388_W_in=> c0_n388_W_in, 
            c0_n389_W_in=> c0_n389_W_in, 
            c0_n390_W_in=> c0_n390_W_in, 
            c0_n391_W_in=> c0_n391_W_in, 
            c0_n392_W_in=> c0_n392_W_in, 
            c0_n393_W_in=> c0_n393_W_in, 
            c0_n394_W_in=> c0_n394_W_in, 
            c0_n395_W_in=> c0_n395_W_in, 
            c0_n396_W_in=> c0_n396_W_in, 
            c0_n397_W_in=> c0_n397_W_in, 
            c0_n398_W_in=> c0_n398_W_in, 
            c0_n399_W_in=> c0_n399_W_in, 
            c0_n400_W_in=> c0_n400_W_in, 
            c0_n401_W_in=> c0_n401_W_in, 
            c0_n402_W_in=> c0_n402_W_in, 
            c0_n403_W_in=> c0_n403_W_in, 
            c0_n404_W_in=> c0_n404_W_in, 
            c0_n405_W_in=> c0_n405_W_in, 
            c0_n406_W_in=> c0_n406_W_in, 
            c0_n407_W_in=> c0_n407_W_in, 
            c0_n408_W_in=> c0_n408_W_in, 
            c0_n409_W_in=> c0_n409_W_in, 
            c0_n410_W_in=> c0_n410_W_in, 
            c0_n411_W_in=> c0_n411_W_in, 
            c0_n412_W_in=> c0_n412_W_in, 
            c0_n413_W_in=> c0_n413_W_in, 
            c0_n414_W_in=> c0_n414_W_in, 
            c0_n415_W_in=> c0_n415_W_in, 
            c0_n416_W_in=> c0_n416_W_in, 
            c0_n417_W_in=> c0_n417_W_in, 
            c0_n418_W_in=> c0_n418_W_in, 
            c0_n419_W_in=> c0_n419_W_in, 
            c0_n420_W_in=> c0_n420_W_in, 
            c0_n421_W_in=> c0_n421_W_in, 
            c0_n422_W_in=> c0_n422_W_in, 
            c0_n423_W_in=> c0_n423_W_in, 
            c0_n424_W_in=> c0_n424_W_in, 
            c0_n425_W_in=> c0_n425_W_in, 
            c0_n426_W_in=> c0_n426_W_in, 
            c0_n427_W_in=> c0_n427_W_in, 
            c0_n428_W_in=> c0_n428_W_in, 
            c0_n429_W_in=> c0_n429_W_in, 
            c0_n430_W_in=> c0_n430_W_in, 
            c0_n431_W_in=> c0_n431_W_in, 
            c0_n432_W_in=> c0_n432_W_in, 
            c0_n433_W_in=> c0_n433_W_in, 
            c0_n434_W_in=> c0_n434_W_in, 
            c0_n435_W_in=> c0_n435_W_in, 
            c0_n436_W_in=> c0_n436_W_in, 
            c0_n437_W_in=> c0_n437_W_in, 
            c0_n438_W_in=> c0_n438_W_in, 
            c0_n439_W_in=> c0_n439_W_in, 
            c0_n440_W_in=> c0_n440_W_in, 
            c0_n441_W_in=> c0_n441_W_in, 
            c0_n442_W_in=> c0_n442_W_in, 
            c0_n443_W_in=> c0_n443_W_in, 
            c0_n444_W_in=> c0_n444_W_in, 
            c0_n445_W_in=> c0_n445_W_in, 
            c0_n446_W_in=> c0_n446_W_in, 
            c0_n447_W_in=> c0_n447_W_in, 
            c0_n448_W_in=> c0_n448_W_in, 
            c0_n449_W_in=> c0_n449_W_in, 
            c0_n450_W_in=> c0_n450_W_in, 
            c0_n451_W_in=> c0_n451_W_in, 
            c0_n452_W_in=> c0_n452_W_in, 
            c0_n453_W_in=> c0_n453_W_in, 
            c0_n454_W_in=> c0_n454_W_in, 
            c0_n455_W_in=> c0_n455_W_in, 
            c0_n456_W_in=> c0_n456_W_in, 
            c0_n457_W_in=> c0_n457_W_in, 
            c0_n458_W_in=> c0_n458_W_in, 
            c0_n459_W_in=> c0_n459_W_in, 
            c0_n460_W_in=> c0_n460_W_in, 
            c0_n461_W_in=> c0_n461_W_in, 
            c0_n462_W_in=> c0_n462_W_in, 
            c0_n463_W_in=> c0_n463_W_in, 
            c0_n464_W_in=> c0_n464_W_in, 
            c0_n465_W_in=> c0_n465_W_in, 
            c0_n466_W_in=> c0_n466_W_in, 
            c0_n467_W_in=> c0_n467_W_in, 
            c0_n468_W_in=> c0_n468_W_in, 
            c0_n469_W_in=> c0_n469_W_in, 
            c0_n470_W_in=> c0_n470_W_in, 
            c0_n471_W_in=> c0_n471_W_in, 
            c0_n472_W_in=> c0_n472_W_in, 
            c0_n473_W_in=> c0_n473_W_in, 
            c0_n474_W_in=> c0_n474_W_in, 
            c0_n475_W_in=> c0_n475_W_in, 
            c0_n476_W_in=> c0_n476_W_in, 
            c0_n477_W_in=> c0_n477_W_in, 
            c0_n478_W_in=> c0_n478_W_in, 
            c0_n479_W_in=> c0_n479_W_in, 
            c0_n480_W_in=> c0_n480_W_in, 
            c0_n481_W_in=> c0_n481_W_in, 
            c0_n482_W_in=> c0_n482_W_in, 
            c0_n483_W_in=> c0_n483_W_in, 
            c0_n484_W_in=> c0_n484_W_in, 
            c0_n485_W_in=> c0_n485_W_in, 
            c0_n486_W_in=> c0_n486_W_in, 
            c0_n487_W_in=> c0_n487_W_in, 
            c0_n488_W_in=> c0_n488_W_in, 
            c0_n489_W_in=> c0_n489_W_in, 
            c0_n490_W_in=> c0_n490_W_in, 
            c0_n491_W_in=> c0_n491_W_in, 
            c0_n492_W_in=> c0_n492_W_in, 
            c0_n493_W_in=> c0_n493_W_in, 
            c0_n494_W_in=> c0_n494_W_in, 
            c0_n495_W_in=> c0_n495_W_in, 
            c0_n496_W_in=> c0_n496_W_in, 
            c0_n497_W_in=> c0_n497_W_in, 
            c0_n498_W_in=> c0_n498_W_in, 
            c0_n499_W_in=> c0_n499_W_in, 
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c0_n0_IO_out=> c0_n0_IO_out, 
            c0_n1_IO_out=> c0_n1_IO_out, 
            c0_n2_IO_out=> c0_n2_IO_out, 
            c0_n3_IO_out=> c0_n3_IO_out, 
            c0_n4_IO_out=> c0_n4_IO_out, 
            c0_n5_IO_out=> c0_n5_IO_out, 
            c0_n6_IO_out=> c0_n6_IO_out, 
            c0_n7_IO_out=> c0_n7_IO_out, 
            c0_n8_IO_out=> c0_n8_IO_out, 
            c0_n9_IO_out=> c0_n9_IO_out, 
            c0_n10_IO_out=> c0_n10_IO_out, 
            c0_n11_IO_out=> c0_n11_IO_out, 
            c0_n12_IO_out=> c0_n12_IO_out, 
            c0_n13_IO_out=> c0_n13_IO_out, 
            c0_n14_IO_out=> c0_n14_IO_out, 
            c0_n15_IO_out=> c0_n15_IO_out, 
            c0_n16_IO_out=> c0_n16_IO_out, 
            c0_n17_IO_out=> c0_n17_IO_out, 
            c0_n18_IO_out=> c0_n18_IO_out, 
            c0_n19_IO_out=> c0_n19_IO_out, 
            c0_n20_IO_out=> c0_n20_IO_out, 
            c0_n21_IO_out=> c0_n21_IO_out, 
            c0_n22_IO_out=> c0_n22_IO_out, 
            c0_n23_IO_out=> c0_n23_IO_out, 
            c0_n24_IO_out=> c0_n24_IO_out, 
            c0_n25_IO_out=> c0_n25_IO_out, 
            c0_n26_IO_out=> c0_n26_IO_out, 
            c0_n27_IO_out=> c0_n27_IO_out, 
            c0_n28_IO_out=> c0_n28_IO_out, 
            c0_n29_IO_out=> c0_n29_IO_out, 
            c0_n30_IO_out=> c0_n30_IO_out, 
            c0_n31_IO_out=> c0_n31_IO_out, 
            c0_n32_IO_out=> c0_n32_IO_out, 
            c0_n33_IO_out=> c0_n33_IO_out, 
            c0_n34_IO_out=> c0_n34_IO_out, 
            c0_n35_IO_out=> c0_n35_IO_out, 
            c0_n36_IO_out=> c0_n36_IO_out, 
            c0_n37_IO_out=> c0_n37_IO_out, 
            c0_n38_IO_out=> c0_n38_IO_out, 
            c0_n39_IO_out=> c0_n39_IO_out, 
            c0_n40_IO_out=> c0_n40_IO_out, 
            c0_n41_IO_out=> c0_n41_IO_out, 
            c0_n42_IO_out=> c0_n42_IO_out, 
            c0_n43_IO_out=> c0_n43_IO_out, 
            c0_n44_IO_out=> c0_n44_IO_out, 
            c0_n45_IO_out=> c0_n45_IO_out, 
            c0_n46_IO_out=> c0_n46_IO_out, 
            c0_n47_IO_out=> c0_n47_IO_out, 
            c0_n48_IO_out=> c0_n48_IO_out, 
            c0_n49_IO_out=> c0_n49_IO_out, 
            c0_n50_IO_out=> c0_n50_IO_out, 
            c0_n51_IO_out=> c0_n51_IO_out, 
            c0_n52_IO_out=> c0_n52_IO_out, 
            c0_n53_IO_out=> c0_n53_IO_out, 
            c0_n54_IO_out=> c0_n54_IO_out, 
            c0_n55_IO_out=> c0_n55_IO_out, 
            c0_n56_IO_out=> c0_n56_IO_out, 
            c0_n57_IO_out=> c0_n57_IO_out, 
            c0_n58_IO_out=> c0_n58_IO_out, 
            c0_n59_IO_out=> c0_n59_IO_out, 
            c0_n60_IO_out=> c0_n60_IO_out, 
            c0_n61_IO_out=> c0_n61_IO_out, 
            c0_n62_IO_out=> c0_n62_IO_out, 
            c0_n63_IO_out=> c0_n63_IO_out, 
            c0_n64_IO_out=> c0_n64_IO_out, 
            c0_n65_IO_out=> c0_n65_IO_out, 
            c0_n66_IO_out=> c0_n66_IO_out, 
            c0_n67_IO_out=> c0_n67_IO_out, 
            c0_n68_IO_out=> c0_n68_IO_out, 
            c0_n69_IO_out=> c0_n69_IO_out, 
            c0_n70_IO_out=> c0_n70_IO_out, 
            c0_n71_IO_out=> c0_n71_IO_out, 
            c0_n72_IO_out=> c0_n72_IO_out, 
            c0_n73_IO_out=> c0_n73_IO_out, 
            c0_n74_IO_out=> c0_n74_IO_out, 
            c0_n75_IO_out=> c0_n75_IO_out, 
            c0_n76_IO_out=> c0_n76_IO_out, 
            c0_n77_IO_out=> c0_n77_IO_out, 
            c0_n78_IO_out=> c0_n78_IO_out, 
            c0_n79_IO_out=> c0_n79_IO_out, 
            c0_n80_IO_out=> c0_n80_IO_out, 
            c0_n81_IO_out=> c0_n81_IO_out, 
            c0_n82_IO_out=> c0_n82_IO_out, 
            c0_n83_IO_out=> c0_n83_IO_out, 
            c0_n84_IO_out=> c0_n84_IO_out, 
            c0_n85_IO_out=> c0_n85_IO_out, 
            c0_n86_IO_out=> c0_n86_IO_out, 
            c0_n87_IO_out=> c0_n87_IO_out, 
            c0_n88_IO_out=> c0_n88_IO_out, 
            c0_n89_IO_out=> c0_n89_IO_out, 
            c0_n90_IO_out=> c0_n90_IO_out, 
            c0_n91_IO_out=> c0_n91_IO_out, 
            c0_n92_IO_out=> c0_n92_IO_out, 
            c0_n93_IO_out=> c0_n93_IO_out, 
            c0_n94_IO_out=> c0_n94_IO_out, 
            c0_n95_IO_out=> c0_n95_IO_out, 
            c0_n96_IO_out=> c0_n96_IO_out, 
            c0_n97_IO_out=> c0_n97_IO_out, 
            c0_n98_IO_out=> c0_n98_IO_out, 
            c0_n99_IO_out=> c0_n99_IO_out, 
            c0_n100_IO_out=> c0_n100_IO_out, 
            c0_n101_IO_out=> c0_n101_IO_out, 
            c0_n102_IO_out=> c0_n102_IO_out, 
            c0_n103_IO_out=> c0_n103_IO_out, 
            c0_n104_IO_out=> c0_n104_IO_out, 
            c0_n105_IO_out=> c0_n105_IO_out, 
            c0_n106_IO_out=> c0_n106_IO_out, 
            c0_n107_IO_out=> c0_n107_IO_out, 
            c0_n108_IO_out=> c0_n108_IO_out, 
            c0_n109_IO_out=> c0_n109_IO_out, 
            c0_n110_IO_out=> c0_n110_IO_out, 
            c0_n111_IO_out=> c0_n111_IO_out, 
            c0_n112_IO_out=> c0_n112_IO_out, 
            c0_n113_IO_out=> c0_n113_IO_out, 
            c0_n114_IO_out=> c0_n114_IO_out, 
            c0_n115_IO_out=> c0_n115_IO_out, 
            c0_n116_IO_out=> c0_n116_IO_out, 
            c0_n117_IO_out=> c0_n117_IO_out, 
            c0_n118_IO_out=> c0_n118_IO_out, 
            c0_n119_IO_out=> c0_n119_IO_out, 
            c0_n120_IO_out=> c0_n120_IO_out, 
            c0_n121_IO_out=> c0_n121_IO_out, 
            c0_n122_IO_out=> c0_n122_IO_out, 
            c0_n123_IO_out=> c0_n123_IO_out, 
            c0_n124_IO_out=> c0_n124_IO_out, 
            c0_n125_IO_out=> c0_n125_IO_out, 
            c0_n126_IO_out=> c0_n126_IO_out, 
            c0_n127_IO_out=> c0_n127_IO_out, 
            c0_n128_IO_out=> c0_n128_IO_out, 
            c0_n129_IO_out=> c0_n129_IO_out, 
            c0_n130_IO_out=> c0_n130_IO_out, 
            c0_n131_IO_out=> c0_n131_IO_out, 
            c0_n132_IO_out=> c0_n132_IO_out, 
            c0_n133_IO_out=> c0_n133_IO_out, 
            c0_n134_IO_out=> c0_n134_IO_out, 
            c0_n135_IO_out=> c0_n135_IO_out, 
            c0_n136_IO_out=> c0_n136_IO_out, 
            c0_n137_IO_out=> c0_n137_IO_out, 
            c0_n138_IO_out=> c0_n138_IO_out, 
            c0_n139_IO_out=> c0_n139_IO_out, 
            c0_n140_IO_out=> c0_n140_IO_out, 
            c0_n141_IO_out=> c0_n141_IO_out, 
            c0_n142_IO_out=> c0_n142_IO_out, 
            c0_n143_IO_out=> c0_n143_IO_out, 
            c0_n144_IO_out=> c0_n144_IO_out, 
            c0_n145_IO_out=> c0_n145_IO_out, 
            c0_n146_IO_out=> c0_n146_IO_out, 
            c0_n147_IO_out=> c0_n147_IO_out, 
            c0_n148_IO_out=> c0_n148_IO_out, 
            c0_n149_IO_out=> c0_n149_IO_out, 
            c0_n150_IO_out=> c0_n150_IO_out, 
            c0_n151_IO_out=> c0_n151_IO_out, 
            c0_n152_IO_out=> c0_n152_IO_out, 
            c0_n153_IO_out=> c0_n153_IO_out, 
            c0_n154_IO_out=> c0_n154_IO_out, 
            c0_n155_IO_out=> c0_n155_IO_out, 
            c0_n156_IO_out=> c0_n156_IO_out, 
            c0_n157_IO_out=> c0_n157_IO_out, 
            c0_n158_IO_out=> c0_n158_IO_out, 
            c0_n159_IO_out=> c0_n159_IO_out, 
            c0_n160_IO_out=> c0_n160_IO_out, 
            c0_n161_IO_out=> c0_n161_IO_out, 
            c0_n162_IO_out=> c0_n162_IO_out, 
            c0_n163_IO_out=> c0_n163_IO_out, 
            c0_n164_IO_out=> c0_n164_IO_out, 
            c0_n165_IO_out=> c0_n165_IO_out, 
            c0_n166_IO_out=> c0_n166_IO_out, 
            c0_n167_IO_out=> c0_n167_IO_out, 
            c0_n168_IO_out=> c0_n168_IO_out, 
            c0_n169_IO_out=> c0_n169_IO_out, 
            c0_n170_IO_out=> c0_n170_IO_out, 
            c0_n171_IO_out=> c0_n171_IO_out, 
            c0_n172_IO_out=> c0_n172_IO_out, 
            c0_n173_IO_out=> c0_n173_IO_out, 
            c0_n174_IO_out=> c0_n174_IO_out, 
            c0_n175_IO_out=> c0_n175_IO_out, 
            c0_n176_IO_out=> c0_n176_IO_out, 
            c0_n177_IO_out=> c0_n177_IO_out, 
            c0_n178_IO_out=> c0_n178_IO_out, 
            c0_n179_IO_out=> c0_n179_IO_out, 
            c0_n180_IO_out=> c0_n180_IO_out, 
            c0_n181_IO_out=> c0_n181_IO_out, 
            c0_n182_IO_out=> c0_n182_IO_out, 
            c0_n183_IO_out=> c0_n183_IO_out, 
            c0_n184_IO_out=> c0_n184_IO_out, 
            c0_n185_IO_out=> c0_n185_IO_out, 
            c0_n186_IO_out=> c0_n186_IO_out, 
            c0_n187_IO_out=> c0_n187_IO_out, 
            c0_n188_IO_out=> c0_n188_IO_out, 
            c0_n189_IO_out=> c0_n189_IO_out, 
            c0_n190_IO_out=> c0_n190_IO_out, 
            c0_n191_IO_out=> c0_n191_IO_out, 
            c0_n192_IO_out=> c0_n192_IO_out, 
            c0_n193_IO_out=> c0_n193_IO_out, 
            c0_n194_IO_out=> c0_n194_IO_out, 
            c0_n195_IO_out=> c0_n195_IO_out, 
            c0_n196_IO_out=> c0_n196_IO_out, 
            c0_n197_IO_out=> c0_n197_IO_out, 
            c0_n198_IO_out=> c0_n198_IO_out, 
            c0_n199_IO_out=> c0_n199_IO_out, 
            c0_n200_IO_out=> c0_n200_IO_out, 
            c0_n201_IO_out=> c0_n201_IO_out, 
            c0_n202_IO_out=> c0_n202_IO_out, 
            c0_n203_IO_out=> c0_n203_IO_out, 
            c0_n204_IO_out=> c0_n204_IO_out, 
            c0_n205_IO_out=> c0_n205_IO_out, 
            c0_n206_IO_out=> c0_n206_IO_out, 
            c0_n207_IO_out=> c0_n207_IO_out, 
            c0_n208_IO_out=> c0_n208_IO_out, 
            c0_n209_IO_out=> c0_n209_IO_out, 
            c0_n210_IO_out=> c0_n210_IO_out, 
            c0_n211_IO_out=> c0_n211_IO_out, 
            c0_n212_IO_out=> c0_n212_IO_out, 
            c0_n213_IO_out=> c0_n213_IO_out, 
            c0_n214_IO_out=> c0_n214_IO_out, 
            c0_n215_IO_out=> c0_n215_IO_out, 
            c0_n216_IO_out=> c0_n216_IO_out, 
            c0_n217_IO_out=> c0_n217_IO_out, 
            c0_n218_IO_out=> c0_n218_IO_out, 
            c0_n219_IO_out=> c0_n219_IO_out, 
            c0_n220_IO_out=> c0_n220_IO_out, 
            c0_n221_IO_out=> c0_n221_IO_out, 
            c0_n222_IO_out=> c0_n222_IO_out, 
            c0_n223_IO_out=> c0_n223_IO_out, 
            c0_n224_IO_out=> c0_n224_IO_out, 
            c0_n225_IO_out=> c0_n225_IO_out, 
            c0_n226_IO_out=> c0_n226_IO_out, 
            c0_n227_IO_out=> c0_n227_IO_out, 
            c0_n228_IO_out=> c0_n228_IO_out, 
            c0_n229_IO_out=> c0_n229_IO_out, 
            c0_n230_IO_out=> c0_n230_IO_out, 
            c0_n231_IO_out=> c0_n231_IO_out, 
            c0_n232_IO_out=> c0_n232_IO_out, 
            c0_n233_IO_out=> c0_n233_IO_out, 
            c0_n234_IO_out=> c0_n234_IO_out, 
            c0_n235_IO_out=> c0_n235_IO_out, 
            c0_n236_IO_out=> c0_n236_IO_out, 
            c0_n237_IO_out=> c0_n237_IO_out, 
            c0_n238_IO_out=> c0_n238_IO_out, 
            c0_n239_IO_out=> c0_n239_IO_out, 
            c0_n240_IO_out=> c0_n240_IO_out, 
            c0_n241_IO_out=> c0_n241_IO_out, 
            c0_n242_IO_out=> c0_n242_IO_out, 
            c0_n243_IO_out=> c0_n243_IO_out, 
            c0_n244_IO_out=> c0_n244_IO_out, 
            c0_n245_IO_out=> c0_n245_IO_out, 
            c0_n246_IO_out=> c0_n246_IO_out, 
            c0_n247_IO_out=> c0_n247_IO_out, 
            c0_n248_IO_out=> c0_n248_IO_out, 
            c0_n249_IO_out=> c0_n249_IO_out, 
            c0_n250_IO_out=> c0_n250_IO_out, 
            c0_n251_IO_out=> c0_n251_IO_out, 
            c0_n252_IO_out=> c0_n252_IO_out, 
            c0_n253_IO_out=> c0_n253_IO_out, 
            c0_n254_IO_out=> c0_n254_IO_out, 
            c0_n255_IO_out=> c0_n255_IO_out, 
            c0_n256_IO_out=> c0_n256_IO_out, 
            c0_n257_IO_out=> c0_n257_IO_out, 
            c0_n258_IO_out=> c0_n258_IO_out, 
            c0_n259_IO_out=> c0_n259_IO_out, 
            c0_n260_IO_out=> c0_n260_IO_out, 
            c0_n261_IO_out=> c0_n261_IO_out, 
            c0_n262_IO_out=> c0_n262_IO_out, 
            c0_n263_IO_out=> c0_n263_IO_out, 
            c0_n264_IO_out=> c0_n264_IO_out, 
            c0_n265_IO_out=> c0_n265_IO_out, 
            c0_n266_IO_out=> c0_n266_IO_out, 
            c0_n267_IO_out=> c0_n267_IO_out, 
            c0_n268_IO_out=> c0_n268_IO_out, 
            c0_n269_IO_out=> c0_n269_IO_out, 
            c0_n270_IO_out=> c0_n270_IO_out, 
            c0_n271_IO_out=> c0_n271_IO_out, 
            c0_n272_IO_out=> c0_n272_IO_out, 
            c0_n273_IO_out=> c0_n273_IO_out, 
            c0_n274_IO_out=> c0_n274_IO_out, 
            c0_n275_IO_out=> c0_n275_IO_out, 
            c0_n276_IO_out=> c0_n276_IO_out, 
            c0_n277_IO_out=> c0_n277_IO_out, 
            c0_n278_IO_out=> c0_n278_IO_out, 
            c0_n279_IO_out=> c0_n279_IO_out, 
            c0_n280_IO_out=> c0_n280_IO_out, 
            c0_n281_IO_out=> c0_n281_IO_out, 
            c0_n282_IO_out=> c0_n282_IO_out, 
            c0_n283_IO_out=> c0_n283_IO_out, 
            c0_n284_IO_out=> c0_n284_IO_out, 
            c0_n285_IO_out=> c0_n285_IO_out, 
            c0_n286_IO_out=> c0_n286_IO_out, 
            c0_n287_IO_out=> c0_n287_IO_out, 
            c0_n288_IO_out=> c0_n288_IO_out, 
            c0_n289_IO_out=> c0_n289_IO_out, 
            c0_n290_IO_out=> c0_n290_IO_out, 
            c0_n291_IO_out=> c0_n291_IO_out, 
            c0_n292_IO_out=> c0_n292_IO_out, 
            c0_n293_IO_out=> c0_n293_IO_out, 
            c0_n294_IO_out=> c0_n294_IO_out, 
            c0_n295_IO_out=> c0_n295_IO_out, 
            c0_n296_IO_out=> c0_n296_IO_out, 
            c0_n297_IO_out=> c0_n297_IO_out, 
            c0_n298_IO_out=> c0_n298_IO_out, 
            c0_n299_IO_out=> c0_n299_IO_out, 
            c0_n300_IO_out=> c0_n300_IO_out, 
            c0_n301_IO_out=> c0_n301_IO_out, 
            c0_n302_IO_out=> c0_n302_IO_out, 
            c0_n303_IO_out=> c0_n303_IO_out, 
            c0_n304_IO_out=> c0_n304_IO_out, 
            c0_n305_IO_out=> c0_n305_IO_out, 
            c0_n306_IO_out=> c0_n306_IO_out, 
            c0_n307_IO_out=> c0_n307_IO_out, 
            c0_n308_IO_out=> c0_n308_IO_out, 
            c0_n309_IO_out=> c0_n309_IO_out, 
            c0_n310_IO_out=> c0_n310_IO_out, 
            c0_n311_IO_out=> c0_n311_IO_out, 
            c0_n312_IO_out=> c0_n312_IO_out, 
            c0_n313_IO_out=> c0_n313_IO_out, 
            c0_n314_IO_out=> c0_n314_IO_out, 
            c0_n315_IO_out=> c0_n315_IO_out, 
            c0_n316_IO_out=> c0_n316_IO_out, 
            c0_n317_IO_out=> c0_n317_IO_out, 
            c0_n318_IO_out=> c0_n318_IO_out, 
            c0_n319_IO_out=> c0_n319_IO_out, 
            c0_n320_IO_out=> c0_n320_IO_out, 
            c0_n321_IO_out=> c0_n321_IO_out, 
            c0_n322_IO_out=> c0_n322_IO_out, 
            c0_n323_IO_out=> c0_n323_IO_out, 
            c0_n324_IO_out=> c0_n324_IO_out, 
            c0_n325_IO_out=> c0_n325_IO_out, 
            c0_n326_IO_out=> c0_n326_IO_out, 
            c0_n327_IO_out=> c0_n327_IO_out, 
            c0_n328_IO_out=> c0_n328_IO_out, 
            c0_n329_IO_out=> c0_n329_IO_out, 
            c0_n330_IO_out=> c0_n330_IO_out, 
            c0_n331_IO_out=> c0_n331_IO_out, 
            c0_n332_IO_out=> c0_n332_IO_out, 
            c0_n333_IO_out=> c0_n333_IO_out, 
            c0_n334_IO_out=> c0_n334_IO_out, 
            c0_n335_IO_out=> c0_n335_IO_out, 
            c0_n336_IO_out=> c0_n336_IO_out, 
            c0_n337_IO_out=> c0_n337_IO_out, 
            c0_n338_IO_out=> c0_n338_IO_out, 
            c0_n339_IO_out=> c0_n339_IO_out, 
            c0_n340_IO_out=> c0_n340_IO_out, 
            c0_n341_IO_out=> c0_n341_IO_out, 
            c0_n342_IO_out=> c0_n342_IO_out, 
            c0_n343_IO_out=> c0_n343_IO_out, 
            c0_n344_IO_out=> c0_n344_IO_out, 
            c0_n345_IO_out=> c0_n345_IO_out, 
            c0_n346_IO_out=> c0_n346_IO_out, 
            c0_n347_IO_out=> c0_n347_IO_out, 
            c0_n348_IO_out=> c0_n348_IO_out, 
            c0_n349_IO_out=> c0_n349_IO_out, 
            c0_n350_IO_out=> c0_n350_IO_out, 
            c0_n351_IO_out=> c0_n351_IO_out, 
            c0_n352_IO_out=> c0_n352_IO_out, 
            c0_n353_IO_out=> c0_n353_IO_out, 
            c0_n354_IO_out=> c0_n354_IO_out, 
            c0_n355_IO_out=> c0_n355_IO_out, 
            c0_n356_IO_out=> c0_n356_IO_out, 
            c0_n357_IO_out=> c0_n357_IO_out, 
            c0_n358_IO_out=> c0_n358_IO_out, 
            c0_n359_IO_out=> c0_n359_IO_out, 
            c0_n360_IO_out=> c0_n360_IO_out, 
            c0_n361_IO_out=> c0_n361_IO_out, 
            c0_n362_IO_out=> c0_n362_IO_out, 
            c0_n363_IO_out=> c0_n363_IO_out, 
            c0_n364_IO_out=> c0_n364_IO_out, 
            c0_n365_IO_out=> c0_n365_IO_out, 
            c0_n366_IO_out=> c0_n366_IO_out, 
            c0_n367_IO_out=> c0_n367_IO_out, 
            c0_n368_IO_out=> c0_n368_IO_out, 
            c0_n369_IO_out=> c0_n369_IO_out, 
            c0_n370_IO_out=> c0_n370_IO_out, 
            c0_n371_IO_out=> c0_n371_IO_out, 
            c0_n372_IO_out=> c0_n372_IO_out, 
            c0_n373_IO_out=> c0_n373_IO_out, 
            c0_n374_IO_out=> c0_n374_IO_out, 
            c0_n375_IO_out=> c0_n375_IO_out, 
            c0_n376_IO_out=> c0_n376_IO_out, 
            c0_n377_IO_out=> c0_n377_IO_out, 
            c0_n378_IO_out=> c0_n378_IO_out, 
            c0_n379_IO_out=> c0_n379_IO_out, 
            c0_n380_IO_out=> c0_n380_IO_out, 
            c0_n381_IO_out=> c0_n381_IO_out, 
            c0_n382_IO_out=> c0_n382_IO_out, 
            c0_n383_IO_out=> c0_n383_IO_out, 
            c0_n384_IO_out=> c0_n384_IO_out, 
            c0_n385_IO_out=> c0_n385_IO_out, 
            c0_n386_IO_out=> c0_n386_IO_out, 
            c0_n387_IO_out=> c0_n387_IO_out, 
            c0_n388_IO_out=> c0_n388_IO_out, 
            c0_n389_IO_out=> c0_n389_IO_out, 
            c0_n390_IO_out=> c0_n390_IO_out, 
            c0_n391_IO_out=> c0_n391_IO_out, 
            c0_n392_IO_out=> c0_n392_IO_out, 
            c0_n393_IO_out=> c0_n393_IO_out, 
            c0_n394_IO_out=> c0_n394_IO_out, 
            c0_n395_IO_out=> c0_n395_IO_out, 
            c0_n396_IO_out=> c0_n396_IO_out, 
            c0_n397_IO_out=> c0_n397_IO_out, 
            c0_n398_IO_out=> c0_n398_IO_out, 
            c0_n399_IO_out=> c0_n399_IO_out, 
            c0_n400_IO_out=> c0_n400_IO_out, 
            c0_n401_IO_out=> c0_n401_IO_out, 
            c0_n402_IO_out=> c0_n402_IO_out, 
            c0_n403_IO_out=> c0_n403_IO_out, 
            c0_n404_IO_out=> c0_n404_IO_out, 
            c0_n405_IO_out=> c0_n405_IO_out, 
            c0_n406_IO_out=> c0_n406_IO_out, 
            c0_n407_IO_out=> c0_n407_IO_out, 
            c0_n408_IO_out=> c0_n408_IO_out, 
            c0_n409_IO_out=> c0_n409_IO_out, 
            c0_n410_IO_out=> c0_n410_IO_out, 
            c0_n411_IO_out=> c0_n411_IO_out, 
            c0_n412_IO_out=> c0_n412_IO_out, 
            c0_n413_IO_out=> c0_n413_IO_out, 
            c0_n414_IO_out=> c0_n414_IO_out, 
            c0_n415_IO_out=> c0_n415_IO_out, 
            c0_n416_IO_out=> c0_n416_IO_out, 
            c0_n417_IO_out=> c0_n417_IO_out, 
            c0_n418_IO_out=> c0_n418_IO_out, 
            c0_n419_IO_out=> c0_n419_IO_out, 
            c0_n420_IO_out=> c0_n420_IO_out, 
            c0_n421_IO_out=> c0_n421_IO_out, 
            c0_n422_IO_out=> c0_n422_IO_out, 
            c0_n423_IO_out=> c0_n423_IO_out, 
            c0_n424_IO_out=> c0_n424_IO_out, 
            c0_n425_IO_out=> c0_n425_IO_out, 
            c0_n426_IO_out=> c0_n426_IO_out, 
            c0_n427_IO_out=> c0_n427_IO_out, 
            c0_n428_IO_out=> c0_n428_IO_out, 
            c0_n429_IO_out=> c0_n429_IO_out, 
            c0_n430_IO_out=> c0_n430_IO_out, 
            c0_n431_IO_out=> c0_n431_IO_out, 
            c0_n432_IO_out=> c0_n432_IO_out, 
            c0_n433_IO_out=> c0_n433_IO_out, 
            c0_n434_IO_out=> c0_n434_IO_out, 
            c0_n435_IO_out=> c0_n435_IO_out, 
            c0_n436_IO_out=> c0_n436_IO_out, 
            c0_n437_IO_out=> c0_n437_IO_out, 
            c0_n438_IO_out=> c0_n438_IO_out, 
            c0_n439_IO_out=> c0_n439_IO_out, 
            c0_n440_IO_out=> c0_n440_IO_out, 
            c0_n441_IO_out=> c0_n441_IO_out, 
            c0_n442_IO_out=> c0_n442_IO_out, 
            c0_n443_IO_out=> c0_n443_IO_out, 
            c0_n444_IO_out=> c0_n444_IO_out, 
            c0_n445_IO_out=> c0_n445_IO_out, 
            c0_n446_IO_out=> c0_n446_IO_out, 
            c0_n447_IO_out=> c0_n447_IO_out, 
            c0_n448_IO_out=> c0_n448_IO_out, 
            c0_n449_IO_out=> c0_n449_IO_out, 
            c0_n450_IO_out=> c0_n450_IO_out, 
            c0_n451_IO_out=> c0_n451_IO_out, 
            c0_n452_IO_out=> c0_n452_IO_out, 
            c0_n453_IO_out=> c0_n453_IO_out, 
            c0_n454_IO_out=> c0_n454_IO_out, 
            c0_n455_IO_out=> c0_n455_IO_out, 
            c0_n456_IO_out=> c0_n456_IO_out, 
            c0_n457_IO_out=> c0_n457_IO_out, 
            c0_n458_IO_out=> c0_n458_IO_out, 
            c0_n459_IO_out=> c0_n459_IO_out, 
            c0_n460_IO_out=> c0_n460_IO_out, 
            c0_n461_IO_out=> c0_n461_IO_out, 
            c0_n462_IO_out=> c0_n462_IO_out, 
            c0_n463_IO_out=> c0_n463_IO_out, 
            c0_n464_IO_out=> c0_n464_IO_out, 
            c0_n465_IO_out=> c0_n465_IO_out, 
            c0_n466_IO_out=> c0_n466_IO_out, 
            c0_n467_IO_out=> c0_n467_IO_out, 
            c0_n468_IO_out=> c0_n468_IO_out, 
            c0_n469_IO_out=> c0_n469_IO_out, 
            c0_n470_IO_out=> c0_n470_IO_out, 
            c0_n471_IO_out=> c0_n471_IO_out, 
            c0_n472_IO_out=> c0_n472_IO_out, 
            c0_n473_IO_out=> c0_n473_IO_out, 
            c0_n474_IO_out=> c0_n474_IO_out, 
            c0_n475_IO_out=> c0_n475_IO_out, 
            c0_n476_IO_out=> c0_n476_IO_out, 
            c0_n477_IO_out=> c0_n477_IO_out, 
            c0_n478_IO_out=> c0_n478_IO_out, 
            c0_n479_IO_out=> c0_n479_IO_out, 
            c0_n480_IO_out=> c0_n480_IO_out, 
            c0_n481_IO_out=> c0_n481_IO_out, 
            c0_n482_IO_out=> c0_n482_IO_out, 
            c0_n483_IO_out=> c0_n483_IO_out, 
            c0_n484_IO_out=> c0_n484_IO_out, 
            c0_n485_IO_out=> c0_n485_IO_out, 
            c0_n486_IO_out=> c0_n486_IO_out, 
            c0_n487_IO_out=> c0_n487_IO_out, 
            c0_n488_IO_out=> c0_n488_IO_out, 
            c0_n489_IO_out=> c0_n489_IO_out, 
            c0_n490_IO_out=> c0_n490_IO_out, 
            c0_n491_IO_out=> c0_n491_IO_out, 
            c0_n492_IO_out=> c0_n492_IO_out, 
            c0_n493_IO_out=> c0_n493_IO_out, 
            c0_n494_IO_out=> c0_n494_IO_out, 
            c0_n495_IO_out=> c0_n495_IO_out, 
            c0_n496_IO_out=> c0_n496_IO_out, 
            c0_n497_IO_out=> c0_n497_IO_out, 
            c0_n498_IO_out=> c0_n498_IO_out, 
            c0_n499_IO_out=> c0_n499_IO_out, 
            -- ['OUT']['manual'] 
            c0_n0_W_out=> c0_n0_W_out, 
            c0_n1_W_out=> c0_n1_W_out, 
            c0_n2_W_out=> c0_n2_W_out, 
            c0_n3_W_out=> c0_n3_W_out, 
            c0_n4_W_out=> c0_n4_W_out, 
            c0_n5_W_out=> c0_n5_W_out, 
            c0_n6_W_out=> c0_n6_W_out, 
            c0_n7_W_out=> c0_n7_W_out, 
            c0_n8_W_out=> c0_n8_W_out, 
            c0_n9_W_out=> c0_n9_W_out, 
            c0_n10_W_out=> c0_n10_W_out, 
            c0_n11_W_out=> c0_n11_W_out, 
            c0_n12_W_out=> c0_n12_W_out, 
            c0_n13_W_out=> c0_n13_W_out, 
            c0_n14_W_out=> c0_n14_W_out, 
            c0_n15_W_out=> c0_n15_W_out, 
            c0_n16_W_out=> c0_n16_W_out, 
            c0_n17_W_out=> c0_n17_W_out, 
            c0_n18_W_out=> c0_n18_W_out, 
            c0_n19_W_out=> c0_n19_W_out, 
            c0_n20_W_out=> c0_n20_W_out, 
            c0_n21_W_out=> c0_n21_W_out, 
            c0_n22_W_out=> c0_n22_W_out, 
            c0_n23_W_out=> c0_n23_W_out, 
            c0_n24_W_out=> c0_n24_W_out, 
            c0_n25_W_out=> c0_n25_W_out, 
            c0_n26_W_out=> c0_n26_W_out, 
            c0_n27_W_out=> c0_n27_W_out, 
            c0_n28_W_out=> c0_n28_W_out, 
            c0_n29_W_out=> c0_n29_W_out, 
            c0_n30_W_out=> c0_n30_W_out, 
            c0_n31_W_out=> c0_n31_W_out, 
            c0_n32_W_out=> c0_n32_W_out, 
            c0_n33_W_out=> c0_n33_W_out, 
            c0_n34_W_out=> c0_n34_W_out, 
            c0_n35_W_out=> c0_n35_W_out, 
            c0_n36_W_out=> c0_n36_W_out, 
            c0_n37_W_out=> c0_n37_W_out, 
            c0_n38_W_out=> c0_n38_W_out, 
            c0_n39_W_out=> c0_n39_W_out, 
            c0_n40_W_out=> c0_n40_W_out, 
            c0_n41_W_out=> c0_n41_W_out, 
            c0_n42_W_out=> c0_n42_W_out, 
            c0_n43_W_out=> c0_n43_W_out, 
            c0_n44_W_out=> c0_n44_W_out, 
            c0_n45_W_out=> c0_n45_W_out, 
            c0_n46_W_out=> c0_n46_W_out, 
            c0_n47_W_out=> c0_n47_W_out, 
            c0_n48_W_out=> c0_n48_W_out, 
            c0_n49_W_out=> c0_n49_W_out, 
            c0_n50_W_out=> c0_n50_W_out, 
            c0_n51_W_out=> c0_n51_W_out, 
            c0_n52_W_out=> c0_n52_W_out, 
            c0_n53_W_out=> c0_n53_W_out, 
            c0_n54_W_out=> c0_n54_W_out, 
            c0_n55_W_out=> c0_n55_W_out, 
            c0_n56_W_out=> c0_n56_W_out, 
            c0_n57_W_out=> c0_n57_W_out, 
            c0_n58_W_out=> c0_n58_W_out, 
            c0_n59_W_out=> c0_n59_W_out, 
            c0_n60_W_out=> c0_n60_W_out, 
            c0_n61_W_out=> c0_n61_W_out, 
            c0_n62_W_out=> c0_n62_W_out, 
            c0_n63_W_out=> c0_n63_W_out, 
            c0_n64_W_out=> c0_n64_W_out, 
            c0_n65_W_out=> c0_n65_W_out, 
            c0_n66_W_out=> c0_n66_W_out, 
            c0_n67_W_out=> c0_n67_W_out, 
            c0_n68_W_out=> c0_n68_W_out, 
            c0_n69_W_out=> c0_n69_W_out, 
            c0_n70_W_out=> c0_n70_W_out, 
            c0_n71_W_out=> c0_n71_W_out, 
            c0_n72_W_out=> c0_n72_W_out, 
            c0_n73_W_out=> c0_n73_W_out, 
            c0_n74_W_out=> c0_n74_W_out, 
            c0_n75_W_out=> c0_n75_W_out, 
            c0_n76_W_out=> c0_n76_W_out, 
            c0_n77_W_out=> c0_n77_W_out, 
            c0_n78_W_out=> c0_n78_W_out, 
            c0_n79_W_out=> c0_n79_W_out, 
            c0_n80_W_out=> c0_n80_W_out, 
            c0_n81_W_out=> c0_n81_W_out, 
            c0_n82_W_out=> c0_n82_W_out, 
            c0_n83_W_out=> c0_n83_W_out, 
            c0_n84_W_out=> c0_n84_W_out, 
            c0_n85_W_out=> c0_n85_W_out, 
            c0_n86_W_out=> c0_n86_W_out, 
            c0_n87_W_out=> c0_n87_W_out, 
            c0_n88_W_out=> c0_n88_W_out, 
            c0_n89_W_out=> c0_n89_W_out, 
            c0_n90_W_out=> c0_n90_W_out, 
            c0_n91_W_out=> c0_n91_W_out, 
            c0_n92_W_out=> c0_n92_W_out, 
            c0_n93_W_out=> c0_n93_W_out, 
            c0_n94_W_out=> c0_n94_W_out, 
            c0_n95_W_out=> c0_n95_W_out, 
            c0_n96_W_out=> c0_n96_W_out, 
            c0_n97_W_out=> c0_n97_W_out, 
            c0_n98_W_out=> c0_n98_W_out, 
            c0_n99_W_out=> c0_n99_W_out, 
            c0_n100_W_out=> c0_n100_W_out, 
            c0_n101_W_out=> c0_n101_W_out, 
            c0_n102_W_out=> c0_n102_W_out, 
            c0_n103_W_out=> c0_n103_W_out, 
            c0_n104_W_out=> c0_n104_W_out, 
            c0_n105_W_out=> c0_n105_W_out, 
            c0_n106_W_out=> c0_n106_W_out, 
            c0_n107_W_out=> c0_n107_W_out, 
            c0_n108_W_out=> c0_n108_W_out, 
            c0_n109_W_out=> c0_n109_W_out, 
            c0_n110_W_out=> c0_n110_W_out, 
            c0_n111_W_out=> c0_n111_W_out, 
            c0_n112_W_out=> c0_n112_W_out, 
            c0_n113_W_out=> c0_n113_W_out, 
            c0_n114_W_out=> c0_n114_W_out, 
            c0_n115_W_out=> c0_n115_W_out, 
            c0_n116_W_out=> c0_n116_W_out, 
            c0_n117_W_out=> c0_n117_W_out, 
            c0_n118_W_out=> c0_n118_W_out, 
            c0_n119_W_out=> c0_n119_W_out, 
            c0_n120_W_out=> c0_n120_W_out, 
            c0_n121_W_out=> c0_n121_W_out, 
            c0_n122_W_out=> c0_n122_W_out, 
            c0_n123_W_out=> c0_n123_W_out, 
            c0_n124_W_out=> c0_n124_W_out, 
            c0_n125_W_out=> c0_n125_W_out, 
            c0_n126_W_out=> c0_n126_W_out, 
            c0_n127_W_out=> c0_n127_W_out, 
            c0_n128_W_out=> c0_n128_W_out, 
            c0_n129_W_out=> c0_n129_W_out, 
            c0_n130_W_out=> c0_n130_W_out, 
            c0_n131_W_out=> c0_n131_W_out, 
            c0_n132_W_out=> c0_n132_W_out, 
            c0_n133_W_out=> c0_n133_W_out, 
            c0_n134_W_out=> c0_n134_W_out, 
            c0_n135_W_out=> c0_n135_W_out, 
            c0_n136_W_out=> c0_n136_W_out, 
            c0_n137_W_out=> c0_n137_W_out, 
            c0_n138_W_out=> c0_n138_W_out, 
            c0_n139_W_out=> c0_n139_W_out, 
            c0_n140_W_out=> c0_n140_W_out, 
            c0_n141_W_out=> c0_n141_W_out, 
            c0_n142_W_out=> c0_n142_W_out, 
            c0_n143_W_out=> c0_n143_W_out, 
            c0_n144_W_out=> c0_n144_W_out, 
            c0_n145_W_out=> c0_n145_W_out, 
            c0_n146_W_out=> c0_n146_W_out, 
            c0_n147_W_out=> c0_n147_W_out, 
            c0_n148_W_out=> c0_n148_W_out, 
            c0_n149_W_out=> c0_n149_W_out, 
            c0_n150_W_out=> c0_n150_W_out, 
            c0_n151_W_out=> c0_n151_W_out, 
            c0_n152_W_out=> c0_n152_W_out, 
            c0_n153_W_out=> c0_n153_W_out, 
            c0_n154_W_out=> c0_n154_W_out, 
            c0_n155_W_out=> c0_n155_W_out, 
            c0_n156_W_out=> c0_n156_W_out, 
            c0_n157_W_out=> c0_n157_W_out, 
            c0_n158_W_out=> c0_n158_W_out, 
            c0_n159_W_out=> c0_n159_W_out, 
            c0_n160_W_out=> c0_n160_W_out, 
            c0_n161_W_out=> c0_n161_W_out, 
            c0_n162_W_out=> c0_n162_W_out, 
            c0_n163_W_out=> c0_n163_W_out, 
            c0_n164_W_out=> c0_n164_W_out, 
            c0_n165_W_out=> c0_n165_W_out, 
            c0_n166_W_out=> c0_n166_W_out, 
            c0_n167_W_out=> c0_n167_W_out, 
            c0_n168_W_out=> c0_n168_W_out, 
            c0_n169_W_out=> c0_n169_W_out, 
            c0_n170_W_out=> c0_n170_W_out, 
            c0_n171_W_out=> c0_n171_W_out, 
            c0_n172_W_out=> c0_n172_W_out, 
            c0_n173_W_out=> c0_n173_W_out, 
            c0_n174_W_out=> c0_n174_W_out, 
            c0_n175_W_out=> c0_n175_W_out, 
            c0_n176_W_out=> c0_n176_W_out, 
            c0_n177_W_out=> c0_n177_W_out, 
            c0_n178_W_out=> c0_n178_W_out, 
            c0_n179_W_out=> c0_n179_W_out, 
            c0_n180_W_out=> c0_n180_W_out, 
            c0_n181_W_out=> c0_n181_W_out, 
            c0_n182_W_out=> c0_n182_W_out, 
            c0_n183_W_out=> c0_n183_W_out, 
            c0_n184_W_out=> c0_n184_W_out, 
            c0_n185_W_out=> c0_n185_W_out, 
            c0_n186_W_out=> c0_n186_W_out, 
            c0_n187_W_out=> c0_n187_W_out, 
            c0_n188_W_out=> c0_n188_W_out, 
            c0_n189_W_out=> c0_n189_W_out, 
            c0_n190_W_out=> c0_n190_W_out, 
            c0_n191_W_out=> c0_n191_W_out, 
            c0_n192_W_out=> c0_n192_W_out, 
            c0_n193_W_out=> c0_n193_W_out, 
            c0_n194_W_out=> c0_n194_W_out, 
            c0_n195_W_out=> c0_n195_W_out, 
            c0_n196_W_out=> c0_n196_W_out, 
            c0_n197_W_out=> c0_n197_W_out, 
            c0_n198_W_out=> c0_n198_W_out, 
            c0_n199_W_out=> c0_n199_W_out, 
            c0_n200_W_out=> c0_n200_W_out, 
            c0_n201_W_out=> c0_n201_W_out, 
            c0_n202_W_out=> c0_n202_W_out, 
            c0_n203_W_out=> c0_n203_W_out, 
            c0_n204_W_out=> c0_n204_W_out, 
            c0_n205_W_out=> c0_n205_W_out, 
            c0_n206_W_out=> c0_n206_W_out, 
            c0_n207_W_out=> c0_n207_W_out, 
            c0_n208_W_out=> c0_n208_W_out, 
            c0_n209_W_out=> c0_n209_W_out, 
            c0_n210_W_out=> c0_n210_W_out, 
            c0_n211_W_out=> c0_n211_W_out, 
            c0_n212_W_out=> c0_n212_W_out, 
            c0_n213_W_out=> c0_n213_W_out, 
            c0_n214_W_out=> c0_n214_W_out, 
            c0_n215_W_out=> c0_n215_W_out, 
            c0_n216_W_out=> c0_n216_W_out, 
            c0_n217_W_out=> c0_n217_W_out, 
            c0_n218_W_out=> c0_n218_W_out, 
            c0_n219_W_out=> c0_n219_W_out, 
            c0_n220_W_out=> c0_n220_W_out, 
            c0_n221_W_out=> c0_n221_W_out, 
            c0_n222_W_out=> c0_n222_W_out, 
            c0_n223_W_out=> c0_n223_W_out, 
            c0_n224_W_out=> c0_n224_W_out, 
            c0_n225_W_out=> c0_n225_W_out, 
            c0_n226_W_out=> c0_n226_W_out, 
            c0_n227_W_out=> c0_n227_W_out, 
            c0_n228_W_out=> c0_n228_W_out, 
            c0_n229_W_out=> c0_n229_W_out, 
            c0_n230_W_out=> c0_n230_W_out, 
            c0_n231_W_out=> c0_n231_W_out, 
            c0_n232_W_out=> c0_n232_W_out, 
            c0_n233_W_out=> c0_n233_W_out, 
            c0_n234_W_out=> c0_n234_W_out, 
            c0_n235_W_out=> c0_n235_W_out, 
            c0_n236_W_out=> c0_n236_W_out, 
            c0_n237_W_out=> c0_n237_W_out, 
            c0_n238_W_out=> c0_n238_W_out, 
            c0_n239_W_out=> c0_n239_W_out, 
            c0_n240_W_out=> c0_n240_W_out, 
            c0_n241_W_out=> c0_n241_W_out, 
            c0_n242_W_out=> c0_n242_W_out, 
            c0_n243_W_out=> c0_n243_W_out, 
            c0_n244_W_out=> c0_n244_W_out, 
            c0_n245_W_out=> c0_n245_W_out, 
            c0_n246_W_out=> c0_n246_W_out, 
            c0_n247_W_out=> c0_n247_W_out, 
            c0_n248_W_out=> c0_n248_W_out, 
            c0_n249_W_out=> c0_n249_W_out, 
            c0_n250_W_out=> c0_n250_W_out, 
            c0_n251_W_out=> c0_n251_W_out, 
            c0_n252_W_out=> c0_n252_W_out, 
            c0_n253_W_out=> c0_n253_W_out, 
            c0_n254_W_out=> c0_n254_W_out, 
            c0_n255_W_out=> c0_n255_W_out, 
            c0_n256_W_out=> c0_n256_W_out, 
            c0_n257_W_out=> c0_n257_W_out, 
            c0_n258_W_out=> c0_n258_W_out, 
            c0_n259_W_out=> c0_n259_W_out, 
            c0_n260_W_out=> c0_n260_W_out, 
            c0_n261_W_out=> c0_n261_W_out, 
            c0_n262_W_out=> c0_n262_W_out, 
            c0_n263_W_out=> c0_n263_W_out, 
            c0_n264_W_out=> c0_n264_W_out, 
            c0_n265_W_out=> c0_n265_W_out, 
            c0_n266_W_out=> c0_n266_W_out, 
            c0_n267_W_out=> c0_n267_W_out, 
            c0_n268_W_out=> c0_n268_W_out, 
            c0_n269_W_out=> c0_n269_W_out, 
            c0_n270_W_out=> c0_n270_W_out, 
            c0_n271_W_out=> c0_n271_W_out, 
            c0_n272_W_out=> c0_n272_W_out, 
            c0_n273_W_out=> c0_n273_W_out, 
            c0_n274_W_out=> c0_n274_W_out, 
            c0_n275_W_out=> c0_n275_W_out, 
            c0_n276_W_out=> c0_n276_W_out, 
            c0_n277_W_out=> c0_n277_W_out, 
            c0_n278_W_out=> c0_n278_W_out, 
            c0_n279_W_out=> c0_n279_W_out, 
            c0_n280_W_out=> c0_n280_W_out, 
            c0_n281_W_out=> c0_n281_W_out, 
            c0_n282_W_out=> c0_n282_W_out, 
            c0_n283_W_out=> c0_n283_W_out, 
            c0_n284_W_out=> c0_n284_W_out, 
            c0_n285_W_out=> c0_n285_W_out, 
            c0_n286_W_out=> c0_n286_W_out, 
            c0_n287_W_out=> c0_n287_W_out, 
            c0_n288_W_out=> c0_n288_W_out, 
            c0_n289_W_out=> c0_n289_W_out, 
            c0_n290_W_out=> c0_n290_W_out, 
            c0_n291_W_out=> c0_n291_W_out, 
            c0_n292_W_out=> c0_n292_W_out, 
            c0_n293_W_out=> c0_n293_W_out, 
            c0_n294_W_out=> c0_n294_W_out, 
            c0_n295_W_out=> c0_n295_W_out, 
            c0_n296_W_out=> c0_n296_W_out, 
            c0_n297_W_out=> c0_n297_W_out, 
            c0_n298_W_out=> c0_n298_W_out, 
            c0_n299_W_out=> c0_n299_W_out, 
            c0_n300_W_out=> c0_n300_W_out, 
            c0_n301_W_out=> c0_n301_W_out, 
            c0_n302_W_out=> c0_n302_W_out, 
            c0_n303_W_out=> c0_n303_W_out, 
            c0_n304_W_out=> c0_n304_W_out, 
            c0_n305_W_out=> c0_n305_W_out, 
            c0_n306_W_out=> c0_n306_W_out, 
            c0_n307_W_out=> c0_n307_W_out, 
            c0_n308_W_out=> c0_n308_W_out, 
            c0_n309_W_out=> c0_n309_W_out, 
            c0_n310_W_out=> c0_n310_W_out, 
            c0_n311_W_out=> c0_n311_W_out, 
            c0_n312_W_out=> c0_n312_W_out, 
            c0_n313_W_out=> c0_n313_W_out, 
            c0_n314_W_out=> c0_n314_W_out, 
            c0_n315_W_out=> c0_n315_W_out, 
            c0_n316_W_out=> c0_n316_W_out, 
            c0_n317_W_out=> c0_n317_W_out, 
            c0_n318_W_out=> c0_n318_W_out, 
            c0_n319_W_out=> c0_n319_W_out, 
            c0_n320_W_out=> c0_n320_W_out, 
            c0_n321_W_out=> c0_n321_W_out, 
            c0_n322_W_out=> c0_n322_W_out, 
            c0_n323_W_out=> c0_n323_W_out, 
            c0_n324_W_out=> c0_n324_W_out, 
            c0_n325_W_out=> c0_n325_W_out, 
            c0_n326_W_out=> c0_n326_W_out, 
            c0_n327_W_out=> c0_n327_W_out, 
            c0_n328_W_out=> c0_n328_W_out, 
            c0_n329_W_out=> c0_n329_W_out, 
            c0_n330_W_out=> c0_n330_W_out, 
            c0_n331_W_out=> c0_n331_W_out, 
            c0_n332_W_out=> c0_n332_W_out, 
            c0_n333_W_out=> c0_n333_W_out, 
            c0_n334_W_out=> c0_n334_W_out, 
            c0_n335_W_out=> c0_n335_W_out, 
            c0_n336_W_out=> c0_n336_W_out, 
            c0_n337_W_out=> c0_n337_W_out, 
            c0_n338_W_out=> c0_n338_W_out, 
            c0_n339_W_out=> c0_n339_W_out, 
            c0_n340_W_out=> c0_n340_W_out, 
            c0_n341_W_out=> c0_n341_W_out, 
            c0_n342_W_out=> c0_n342_W_out, 
            c0_n343_W_out=> c0_n343_W_out, 
            c0_n344_W_out=> c0_n344_W_out, 
            c0_n345_W_out=> c0_n345_W_out, 
            c0_n346_W_out=> c0_n346_W_out, 
            c0_n347_W_out=> c0_n347_W_out, 
            c0_n348_W_out=> c0_n348_W_out, 
            c0_n349_W_out=> c0_n349_W_out, 
            c0_n350_W_out=> c0_n350_W_out, 
            c0_n351_W_out=> c0_n351_W_out, 
            c0_n352_W_out=> c0_n352_W_out, 
            c0_n353_W_out=> c0_n353_W_out, 
            c0_n354_W_out=> c0_n354_W_out, 
            c0_n355_W_out=> c0_n355_W_out, 
            c0_n356_W_out=> c0_n356_W_out, 
            c0_n357_W_out=> c0_n357_W_out, 
            c0_n358_W_out=> c0_n358_W_out, 
            c0_n359_W_out=> c0_n359_W_out, 
            c0_n360_W_out=> c0_n360_W_out, 
            c0_n361_W_out=> c0_n361_W_out, 
            c0_n362_W_out=> c0_n362_W_out, 
            c0_n363_W_out=> c0_n363_W_out, 
            c0_n364_W_out=> c0_n364_W_out, 
            c0_n365_W_out=> c0_n365_W_out, 
            c0_n366_W_out=> c0_n366_W_out, 
            c0_n367_W_out=> c0_n367_W_out, 
            c0_n368_W_out=> c0_n368_W_out, 
            c0_n369_W_out=> c0_n369_W_out, 
            c0_n370_W_out=> c0_n370_W_out, 
            c0_n371_W_out=> c0_n371_W_out, 
            c0_n372_W_out=> c0_n372_W_out, 
            c0_n373_W_out=> c0_n373_W_out, 
            c0_n374_W_out=> c0_n374_W_out, 
            c0_n375_W_out=> c0_n375_W_out, 
            c0_n376_W_out=> c0_n376_W_out, 
            c0_n377_W_out=> c0_n377_W_out, 
            c0_n378_W_out=> c0_n378_W_out, 
            c0_n379_W_out=> c0_n379_W_out, 
            c0_n380_W_out=> c0_n380_W_out, 
            c0_n381_W_out=> c0_n381_W_out, 
            c0_n382_W_out=> c0_n382_W_out, 
            c0_n383_W_out=> c0_n383_W_out, 
            c0_n384_W_out=> c0_n384_W_out, 
            c0_n385_W_out=> c0_n385_W_out, 
            c0_n386_W_out=> c0_n386_W_out, 
            c0_n387_W_out=> c0_n387_W_out, 
            c0_n388_W_out=> c0_n388_W_out, 
            c0_n389_W_out=> c0_n389_W_out, 
            c0_n390_W_out=> c0_n390_W_out, 
            c0_n391_W_out=> c0_n391_W_out, 
            c0_n392_W_out=> c0_n392_W_out, 
            c0_n393_W_out=> c0_n393_W_out, 
            c0_n394_W_out=> c0_n394_W_out, 
            c0_n395_W_out=> c0_n395_W_out, 
            c0_n396_W_out=> c0_n396_W_out, 
            c0_n397_W_out=> c0_n397_W_out, 
            c0_n398_W_out=> c0_n398_W_out, 
            c0_n399_W_out=> c0_n399_W_out, 
            c0_n400_W_out=> c0_n400_W_out, 
            c0_n401_W_out=> c0_n401_W_out, 
            c0_n402_W_out=> c0_n402_W_out, 
            c0_n403_W_out=> c0_n403_W_out, 
            c0_n404_W_out=> c0_n404_W_out, 
            c0_n405_W_out=> c0_n405_W_out, 
            c0_n406_W_out=> c0_n406_W_out, 
            c0_n407_W_out=> c0_n407_W_out, 
            c0_n408_W_out=> c0_n408_W_out, 
            c0_n409_W_out=> c0_n409_W_out, 
            c0_n410_W_out=> c0_n410_W_out, 
            c0_n411_W_out=> c0_n411_W_out, 
            c0_n412_W_out=> c0_n412_W_out, 
            c0_n413_W_out=> c0_n413_W_out, 
            c0_n414_W_out=> c0_n414_W_out, 
            c0_n415_W_out=> c0_n415_W_out, 
            c0_n416_W_out=> c0_n416_W_out, 
            c0_n417_W_out=> c0_n417_W_out, 
            c0_n418_W_out=> c0_n418_W_out, 
            c0_n419_W_out=> c0_n419_W_out, 
            c0_n420_W_out=> c0_n420_W_out, 
            c0_n421_W_out=> c0_n421_W_out, 
            c0_n422_W_out=> c0_n422_W_out, 
            c0_n423_W_out=> c0_n423_W_out, 
            c0_n424_W_out=> c0_n424_W_out, 
            c0_n425_W_out=> c0_n425_W_out, 
            c0_n426_W_out=> c0_n426_W_out, 
            c0_n427_W_out=> c0_n427_W_out, 
            c0_n428_W_out=> c0_n428_W_out, 
            c0_n429_W_out=> c0_n429_W_out, 
            c0_n430_W_out=> c0_n430_W_out, 
            c0_n431_W_out=> c0_n431_W_out, 
            c0_n432_W_out=> c0_n432_W_out, 
            c0_n433_W_out=> c0_n433_W_out, 
            c0_n434_W_out=> c0_n434_W_out, 
            c0_n435_W_out=> c0_n435_W_out, 
            c0_n436_W_out=> c0_n436_W_out, 
            c0_n437_W_out=> c0_n437_W_out, 
            c0_n438_W_out=> c0_n438_W_out, 
            c0_n439_W_out=> c0_n439_W_out, 
            c0_n440_W_out=> c0_n440_W_out, 
            c0_n441_W_out=> c0_n441_W_out, 
            c0_n442_W_out=> c0_n442_W_out, 
            c0_n443_W_out=> c0_n443_W_out, 
            c0_n444_W_out=> c0_n444_W_out, 
            c0_n445_W_out=> c0_n445_W_out, 
            c0_n446_W_out=> c0_n446_W_out, 
            c0_n447_W_out=> c0_n447_W_out, 
            c0_n448_W_out=> c0_n448_W_out, 
            c0_n449_W_out=> c0_n449_W_out, 
            c0_n450_W_out=> c0_n450_W_out, 
            c0_n451_W_out=> c0_n451_W_out, 
            c0_n452_W_out=> c0_n452_W_out, 
            c0_n453_W_out=> c0_n453_W_out, 
            c0_n454_W_out=> c0_n454_W_out, 
            c0_n455_W_out=> c0_n455_W_out, 
            c0_n456_W_out=> c0_n456_W_out, 
            c0_n457_W_out=> c0_n457_W_out, 
            c0_n458_W_out=> c0_n458_W_out, 
            c0_n459_W_out=> c0_n459_W_out, 
            c0_n460_W_out=> c0_n460_W_out, 
            c0_n461_W_out=> c0_n461_W_out, 
            c0_n462_W_out=> c0_n462_W_out, 
            c0_n463_W_out=> c0_n463_W_out, 
            c0_n464_W_out=> c0_n464_W_out, 
            c0_n465_W_out=> c0_n465_W_out, 
            c0_n466_W_out=> c0_n466_W_out, 
            c0_n467_W_out=> c0_n467_W_out, 
            c0_n468_W_out=> c0_n468_W_out, 
            c0_n469_W_out=> c0_n469_W_out, 
            c0_n470_W_out=> c0_n470_W_out, 
            c0_n471_W_out=> c0_n471_W_out, 
            c0_n472_W_out=> c0_n472_W_out, 
            c0_n473_W_out=> c0_n473_W_out, 
            c0_n474_W_out=> c0_n474_W_out, 
            c0_n475_W_out=> c0_n475_W_out, 
            c0_n476_W_out=> c0_n476_W_out, 
            c0_n477_W_out=> c0_n477_W_out, 
            c0_n478_W_out=> c0_n478_W_out, 
            c0_n479_W_out=> c0_n479_W_out, 
            c0_n480_W_out=> c0_n480_W_out, 
            c0_n481_W_out=> c0_n481_W_out, 
            c0_n482_W_out=> c0_n482_W_out, 
            c0_n483_W_out=> c0_n483_W_out, 
            c0_n484_W_out=> c0_n484_W_out, 
            c0_n485_W_out=> c0_n485_W_out, 
            c0_n486_W_out=> c0_n486_W_out, 
            c0_n487_W_out=> c0_n487_W_out, 
            c0_n488_W_out=> c0_n488_W_out, 
            c0_n489_W_out=> c0_n489_W_out, 
            c0_n490_W_out=> c0_n490_W_out, 
            c0_n491_W_out=> c0_n491_W_out, 
            c0_n492_W_out=> c0_n492_W_out, 
            c0_n493_W_out=> c0_n493_W_out, 
            c0_n494_W_out=> c0_n494_W_out, 
            c0_n495_W_out=> c0_n495_W_out, 
            c0_n496_W_out=> c0_n496_W_out, 
            c0_n497_W_out=> c0_n497_W_out, 
            c0_n498_W_out=> c0_n498_W_out, 
            c0_n499_W_out=> c0_n499_W_out
   );
            
camada1_inst_1: ENTITY work.camada1_ReLU_300neuron_8bits_500n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c1_IO_in, 
            c1_n0_W_in=> c0_n0_W_out,
            c1_n1_W_in=> c0_n1_W_out,
            c1_n2_W_in=> c0_n2_W_out,
            c1_n3_W_in=> c0_n3_W_out,
            c1_n4_W_in=> c0_n4_W_out,
            c1_n5_W_in=> c0_n5_W_out,
            c1_n6_W_in=> c0_n6_W_out,
            c1_n7_W_in=> c0_n7_W_out,
            c1_n8_W_in=> c0_n8_W_out,
            c1_n9_W_in=> c0_n9_W_out,
            c1_n10_W_in=> c0_n10_W_out,
            c1_n11_W_in=> c0_n11_W_out,
            c1_n12_W_in=> c0_n12_W_out,
            c1_n13_W_in=> c0_n13_W_out,
            c1_n14_W_in=> c0_n14_W_out,
            c1_n15_W_in=> c0_n15_W_out,
            c1_n16_W_in=> c0_n16_W_out,
            c1_n17_W_in=> c0_n17_W_out,
            c1_n18_W_in=> c0_n18_W_out,
            c1_n19_W_in=> c0_n19_W_out,
            c1_n20_W_in=> c0_n20_W_out,
            c1_n21_W_in=> c0_n21_W_out,
            c1_n22_W_in=> c0_n22_W_out,
            c1_n23_W_in=> c0_n23_W_out,
            c1_n24_W_in=> c0_n24_W_out,
            c1_n25_W_in=> c0_n25_W_out,
            c1_n26_W_in=> c0_n26_W_out,
            c1_n27_W_in=> c0_n27_W_out,
            c1_n28_W_in=> c0_n28_W_out,
            c1_n29_W_in=> c0_n29_W_out,
            c1_n30_W_in=> c0_n30_W_out,
            c1_n31_W_in=> c0_n31_W_out,
            c1_n32_W_in=> c0_n32_W_out,
            c1_n33_W_in=> c0_n33_W_out,
            c1_n34_W_in=> c0_n34_W_out,
            c1_n35_W_in=> c0_n35_W_out,
            c1_n36_W_in=> c0_n36_W_out,
            c1_n37_W_in=> c0_n37_W_out,
            c1_n38_W_in=> c0_n38_W_out,
            c1_n39_W_in=> c0_n39_W_out,
            c1_n40_W_in=> c0_n40_W_out,
            c1_n41_W_in=> c0_n41_W_out,
            c1_n42_W_in=> c0_n42_W_out,
            c1_n43_W_in=> c0_n43_W_out,
            c1_n44_W_in=> c0_n44_W_out,
            c1_n45_W_in=> c0_n45_W_out,
            c1_n46_W_in=> c0_n46_W_out,
            c1_n47_W_in=> c0_n47_W_out,
            c1_n48_W_in=> c0_n48_W_out,
            c1_n49_W_in=> c0_n49_W_out,
            c1_n50_W_in=> c0_n50_W_out,
            c1_n51_W_in=> c0_n51_W_out,
            c1_n52_W_in=> c0_n52_W_out,
            c1_n53_W_in=> c0_n53_W_out,
            c1_n54_W_in=> c0_n54_W_out,
            c1_n55_W_in=> c0_n55_W_out,
            c1_n56_W_in=> c0_n56_W_out,
            c1_n57_W_in=> c0_n57_W_out,
            c1_n58_W_in=> c0_n58_W_out,
            c1_n59_W_in=> c0_n59_W_out,
            c1_n60_W_in=> c0_n60_W_out,
            c1_n61_W_in=> c0_n61_W_out,
            c1_n62_W_in=> c0_n62_W_out,
            c1_n63_W_in=> c0_n63_W_out,
            c1_n64_W_in=> c0_n64_W_out,
            c1_n65_W_in=> c0_n65_W_out,
            c1_n66_W_in=> c0_n66_W_out,
            c1_n67_W_in=> c0_n67_W_out,
            c1_n68_W_in=> c0_n68_W_out,
            c1_n69_W_in=> c0_n69_W_out,
            c1_n70_W_in=> c0_n70_W_out,
            c1_n71_W_in=> c0_n71_W_out,
            c1_n72_W_in=> c0_n72_W_out,
            c1_n73_W_in=> c0_n73_W_out,
            c1_n74_W_in=> c0_n74_W_out,
            c1_n75_W_in=> c0_n75_W_out,
            c1_n76_W_in=> c0_n76_W_out,
            c1_n77_W_in=> c0_n77_W_out,
            c1_n78_W_in=> c0_n78_W_out,
            c1_n79_W_in=> c0_n79_W_out,
            c1_n80_W_in=> c0_n80_W_out,
            c1_n81_W_in=> c0_n81_W_out,
            c1_n82_W_in=> c0_n82_W_out,
            c1_n83_W_in=> c0_n83_W_out,
            c1_n84_W_in=> c0_n84_W_out,
            c1_n85_W_in=> c0_n85_W_out,
            c1_n86_W_in=> c0_n86_W_out,
            c1_n87_W_in=> c0_n87_W_out,
            c1_n88_W_in=> c0_n88_W_out,
            c1_n89_W_in=> c0_n89_W_out,
            c1_n90_W_in=> c0_n90_W_out,
            c1_n91_W_in=> c0_n91_W_out,
            c1_n92_W_in=> c0_n92_W_out,
            c1_n93_W_in=> c0_n93_W_out,
            c1_n94_W_in=> c0_n94_W_out,
            c1_n95_W_in=> c0_n95_W_out,
            c1_n96_W_in=> c0_n96_W_out,
            c1_n97_W_in=> c0_n97_W_out,
            c1_n98_W_in=> c0_n98_W_out,
            c1_n99_W_in=> c0_n99_W_out,
            c1_n100_W_in=> c0_n100_W_out,
            c1_n101_W_in=> c0_n101_W_out,
            c1_n102_W_in=> c0_n102_W_out,
            c1_n103_W_in=> c0_n103_W_out,
            c1_n104_W_in=> c0_n104_W_out,
            c1_n105_W_in=> c0_n105_W_out,
            c1_n106_W_in=> c0_n106_W_out,
            c1_n107_W_in=> c0_n107_W_out,
            c1_n108_W_in=> c0_n108_W_out,
            c1_n109_W_in=> c0_n109_W_out,
            c1_n110_W_in=> c0_n110_W_out,
            c1_n111_W_in=> c0_n111_W_out,
            c1_n112_W_in=> c0_n112_W_out,
            c1_n113_W_in=> c0_n113_W_out,
            c1_n114_W_in=> c0_n114_W_out,
            c1_n115_W_in=> c0_n115_W_out,
            c1_n116_W_in=> c0_n116_W_out,
            c1_n117_W_in=> c0_n117_W_out,
            c1_n118_W_in=> c0_n118_W_out,
            c1_n119_W_in=> c0_n119_W_out,
            c1_n120_W_in=> c0_n120_W_out,
            c1_n121_W_in=> c0_n121_W_out,
            c1_n122_W_in=> c0_n122_W_out,
            c1_n123_W_in=> c0_n123_W_out,
            c1_n124_W_in=> c0_n124_W_out,
            c1_n125_W_in=> c0_n125_W_out,
            c1_n126_W_in=> c0_n126_W_out,
            c1_n127_W_in=> c0_n127_W_out,
            c1_n128_W_in=> c0_n128_W_out,
            c1_n129_W_in=> c0_n129_W_out,
            c1_n130_W_in=> c0_n130_W_out,
            c1_n131_W_in=> c0_n131_W_out,
            c1_n132_W_in=> c0_n132_W_out,
            c1_n133_W_in=> c0_n133_W_out,
            c1_n134_W_in=> c0_n134_W_out,
            c1_n135_W_in=> c0_n135_W_out,
            c1_n136_W_in=> c0_n136_W_out,
            c1_n137_W_in=> c0_n137_W_out,
            c1_n138_W_in=> c0_n138_W_out,
            c1_n139_W_in=> c0_n139_W_out,
            c1_n140_W_in=> c0_n140_W_out,
            c1_n141_W_in=> c0_n141_W_out,
            c1_n142_W_in=> c0_n142_W_out,
            c1_n143_W_in=> c0_n143_W_out,
            c1_n144_W_in=> c0_n144_W_out,
            c1_n145_W_in=> c0_n145_W_out,
            c1_n146_W_in=> c0_n146_W_out,
            c1_n147_W_in=> c0_n147_W_out,
            c1_n148_W_in=> c0_n148_W_out,
            c1_n149_W_in=> c0_n149_W_out,
            c1_n150_W_in=> c0_n150_W_out,
            c1_n151_W_in=> c0_n151_W_out,
            c1_n152_W_in=> c0_n152_W_out,
            c1_n153_W_in=> c0_n153_W_out,
            c1_n154_W_in=> c0_n154_W_out,
            c1_n155_W_in=> c0_n155_W_out,
            c1_n156_W_in=> c0_n156_W_out,
            c1_n157_W_in=> c0_n157_W_out,
            c1_n158_W_in=> c0_n158_W_out,
            c1_n159_W_in=> c0_n159_W_out,
            c1_n160_W_in=> c0_n160_W_out,
            c1_n161_W_in=> c0_n161_W_out,
            c1_n162_W_in=> c0_n162_W_out,
            c1_n163_W_in=> c0_n163_W_out,
            c1_n164_W_in=> c0_n164_W_out,
            c1_n165_W_in=> c0_n165_W_out,
            c1_n166_W_in=> c0_n166_W_out,
            c1_n167_W_in=> c0_n167_W_out,
            c1_n168_W_in=> c0_n168_W_out,
            c1_n169_W_in=> c0_n169_W_out,
            c1_n170_W_in=> c0_n170_W_out,
            c1_n171_W_in=> c0_n171_W_out,
            c1_n172_W_in=> c0_n172_W_out,
            c1_n173_W_in=> c0_n173_W_out,
            c1_n174_W_in=> c0_n174_W_out,
            c1_n175_W_in=> c0_n175_W_out,
            c1_n176_W_in=> c0_n176_W_out,
            c1_n177_W_in=> c0_n177_W_out,
            c1_n178_W_in=> c0_n178_W_out,
            c1_n179_W_in=> c0_n179_W_out,
            c1_n180_W_in=> c0_n180_W_out,
            c1_n181_W_in=> c0_n181_W_out,
            c1_n182_W_in=> c0_n182_W_out,
            c1_n183_W_in=> c0_n183_W_out,
            c1_n184_W_in=> c0_n184_W_out,
            c1_n185_W_in=> c0_n185_W_out,
            c1_n186_W_in=> c0_n186_W_out,
            c1_n187_W_in=> c0_n187_W_out,
            c1_n188_W_in=> c0_n188_W_out,
            c1_n189_W_in=> c0_n189_W_out,
            c1_n190_W_in=> c0_n190_W_out,
            c1_n191_W_in=> c0_n191_W_out,
            c1_n192_W_in=> c0_n192_W_out,
            c1_n193_W_in=> c0_n193_W_out,
            c1_n194_W_in=> c0_n194_W_out,
            c1_n195_W_in=> c0_n195_W_out,
            c1_n196_W_in=> c0_n196_W_out,
            c1_n197_W_in=> c0_n197_W_out,
            c1_n198_W_in=> c0_n198_W_out,
            c1_n199_W_in=> c0_n199_W_out,
            c1_n200_W_in=> c0_n200_W_out,
            c1_n201_W_in=> c0_n201_W_out,
            c1_n202_W_in=> c0_n202_W_out,
            c1_n203_W_in=> c0_n203_W_out,
            c1_n204_W_in=> c0_n204_W_out,
            c1_n205_W_in=> c0_n205_W_out,
            c1_n206_W_in=> c0_n206_W_out,
            c1_n207_W_in=> c0_n207_W_out,
            c1_n208_W_in=> c0_n208_W_out,
            c1_n209_W_in=> c0_n209_W_out,
            c1_n210_W_in=> c0_n210_W_out,
            c1_n211_W_in=> c0_n211_W_out,
            c1_n212_W_in=> c0_n212_W_out,
            c1_n213_W_in=> c0_n213_W_out,
            c1_n214_W_in=> c0_n214_W_out,
            c1_n215_W_in=> c0_n215_W_out,
            c1_n216_W_in=> c0_n216_W_out,
            c1_n217_W_in=> c0_n217_W_out,
            c1_n218_W_in=> c0_n218_W_out,
            c1_n219_W_in=> c0_n219_W_out,
            c1_n220_W_in=> c0_n220_W_out,
            c1_n221_W_in=> c0_n221_W_out,
            c1_n222_W_in=> c0_n222_W_out,
            c1_n223_W_in=> c0_n223_W_out,
            c1_n224_W_in=> c0_n224_W_out,
            c1_n225_W_in=> c0_n225_W_out,
            c1_n226_W_in=> c0_n226_W_out,
            c1_n227_W_in=> c0_n227_W_out,
            c1_n228_W_in=> c0_n228_W_out,
            c1_n229_W_in=> c0_n229_W_out,
            c1_n230_W_in=> c0_n230_W_out,
            c1_n231_W_in=> c0_n231_W_out,
            c1_n232_W_in=> c0_n232_W_out,
            c1_n233_W_in=> c0_n233_W_out,
            c1_n234_W_in=> c0_n234_W_out,
            c1_n235_W_in=> c0_n235_W_out,
            c1_n236_W_in=> c0_n236_W_out,
            c1_n237_W_in=> c0_n237_W_out,
            c1_n238_W_in=> c0_n238_W_out,
            c1_n239_W_in=> c0_n239_W_out,
            c1_n240_W_in=> c0_n240_W_out,
            c1_n241_W_in=> c0_n241_W_out,
            c1_n242_W_in=> c0_n242_W_out,
            c1_n243_W_in=> c0_n243_W_out,
            c1_n244_W_in=> c0_n244_W_out,
            c1_n245_W_in=> c0_n245_W_out,
            c1_n246_W_in=> c0_n246_W_out,
            c1_n247_W_in=> c0_n247_W_out,
            c1_n248_W_in=> c0_n248_W_out,
            c1_n249_W_in=> c0_n249_W_out,
            c1_n250_W_in=> c0_n250_W_out,
            c1_n251_W_in=> c0_n251_W_out,
            c1_n252_W_in=> c0_n252_W_out,
            c1_n253_W_in=> c0_n253_W_out,
            c1_n254_W_in=> c0_n254_W_out,
            c1_n255_W_in=> c0_n255_W_out,
            c1_n256_W_in=> c0_n256_W_out,
            c1_n257_W_in=> c0_n257_W_out,
            c1_n258_W_in=> c0_n258_W_out,
            c1_n259_W_in=> c0_n259_W_out,
            c1_n260_W_in=> c0_n260_W_out,
            c1_n261_W_in=> c0_n261_W_out,
            c1_n262_W_in=> c0_n262_W_out,
            c1_n263_W_in=> c0_n263_W_out,
            c1_n264_W_in=> c0_n264_W_out,
            c1_n265_W_in=> c0_n265_W_out,
            c1_n266_W_in=> c0_n266_W_out,
            c1_n267_W_in=> c0_n267_W_out,
            c1_n268_W_in=> c0_n268_W_out,
            c1_n269_W_in=> c0_n269_W_out,
            c1_n270_W_in=> c0_n270_W_out,
            c1_n271_W_in=> c0_n271_W_out,
            c1_n272_W_in=> c0_n272_W_out,
            c1_n273_W_in=> c0_n273_W_out,
            c1_n274_W_in=> c0_n274_W_out,
            c1_n275_W_in=> c0_n275_W_out,
            c1_n276_W_in=> c0_n276_W_out,
            c1_n277_W_in=> c0_n277_W_out,
            c1_n278_W_in=> c0_n278_W_out,
            c1_n279_W_in=> c0_n279_W_out,
            c1_n280_W_in=> c0_n280_W_out,
            c1_n281_W_in=> c0_n281_W_out,
            c1_n282_W_in=> c0_n282_W_out,
            c1_n283_W_in=> c0_n283_W_out,
            c1_n284_W_in=> c0_n284_W_out,
            c1_n285_W_in=> c0_n285_W_out,
            c1_n286_W_in=> c0_n286_W_out,
            c1_n287_W_in=> c0_n287_W_out,
            c1_n288_W_in=> c0_n288_W_out,
            c1_n289_W_in=> c0_n289_W_out,
            c1_n290_W_in=> c0_n290_W_out,
            c1_n291_W_in=> c0_n291_W_out,
            c1_n292_W_in=> c0_n292_W_out,
            c1_n293_W_in=> c0_n293_W_out,
            c1_n294_W_in=> c0_n294_W_out,
            c1_n295_W_in=> c0_n295_W_out,
            c1_n296_W_in=> c0_n296_W_out,
            c1_n297_W_in=> c0_n297_W_out,
            c1_n298_W_in=> c0_n298_W_out,
            c1_n299_W_in=> c0_n299_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c1_n0_IO_out=> c1_n0_IO_out, 
            c1_n1_IO_out=> c1_n1_IO_out, 
            c1_n2_IO_out=> c1_n2_IO_out, 
            c1_n3_IO_out=> c1_n3_IO_out, 
            c1_n4_IO_out=> c1_n4_IO_out, 
            c1_n5_IO_out=> c1_n5_IO_out, 
            c1_n6_IO_out=> c1_n6_IO_out, 
            c1_n7_IO_out=> c1_n7_IO_out, 
            c1_n8_IO_out=> c1_n8_IO_out, 
            c1_n9_IO_out=> c1_n9_IO_out, 
            c1_n10_IO_out=> c1_n10_IO_out, 
            c1_n11_IO_out=> c1_n11_IO_out, 
            c1_n12_IO_out=> c1_n12_IO_out, 
            c1_n13_IO_out=> c1_n13_IO_out, 
            c1_n14_IO_out=> c1_n14_IO_out, 
            c1_n15_IO_out=> c1_n15_IO_out, 
            c1_n16_IO_out=> c1_n16_IO_out, 
            c1_n17_IO_out=> c1_n17_IO_out, 
            c1_n18_IO_out=> c1_n18_IO_out, 
            c1_n19_IO_out=> c1_n19_IO_out, 
            c1_n20_IO_out=> c1_n20_IO_out, 
            c1_n21_IO_out=> c1_n21_IO_out, 
            c1_n22_IO_out=> c1_n22_IO_out, 
            c1_n23_IO_out=> c1_n23_IO_out, 
            c1_n24_IO_out=> c1_n24_IO_out, 
            c1_n25_IO_out=> c1_n25_IO_out, 
            c1_n26_IO_out=> c1_n26_IO_out, 
            c1_n27_IO_out=> c1_n27_IO_out, 
            c1_n28_IO_out=> c1_n28_IO_out, 
            c1_n29_IO_out=> c1_n29_IO_out, 
            c1_n30_IO_out=> c1_n30_IO_out, 
            c1_n31_IO_out=> c1_n31_IO_out, 
            c1_n32_IO_out=> c1_n32_IO_out, 
            c1_n33_IO_out=> c1_n33_IO_out, 
            c1_n34_IO_out=> c1_n34_IO_out, 
            c1_n35_IO_out=> c1_n35_IO_out, 
            c1_n36_IO_out=> c1_n36_IO_out, 
            c1_n37_IO_out=> c1_n37_IO_out, 
            c1_n38_IO_out=> c1_n38_IO_out, 
            c1_n39_IO_out=> c1_n39_IO_out, 
            c1_n40_IO_out=> c1_n40_IO_out, 
            c1_n41_IO_out=> c1_n41_IO_out, 
            c1_n42_IO_out=> c1_n42_IO_out, 
            c1_n43_IO_out=> c1_n43_IO_out, 
            c1_n44_IO_out=> c1_n44_IO_out, 
            c1_n45_IO_out=> c1_n45_IO_out, 
            c1_n46_IO_out=> c1_n46_IO_out, 
            c1_n47_IO_out=> c1_n47_IO_out, 
            c1_n48_IO_out=> c1_n48_IO_out, 
            c1_n49_IO_out=> c1_n49_IO_out, 
            c1_n50_IO_out=> c1_n50_IO_out, 
            c1_n51_IO_out=> c1_n51_IO_out, 
            c1_n52_IO_out=> c1_n52_IO_out, 
            c1_n53_IO_out=> c1_n53_IO_out, 
            c1_n54_IO_out=> c1_n54_IO_out, 
            c1_n55_IO_out=> c1_n55_IO_out, 
            c1_n56_IO_out=> c1_n56_IO_out, 
            c1_n57_IO_out=> c1_n57_IO_out, 
            c1_n58_IO_out=> c1_n58_IO_out, 
            c1_n59_IO_out=> c1_n59_IO_out, 
            c1_n60_IO_out=> c1_n60_IO_out, 
            c1_n61_IO_out=> c1_n61_IO_out, 
            c1_n62_IO_out=> c1_n62_IO_out, 
            c1_n63_IO_out=> c1_n63_IO_out, 
            c1_n64_IO_out=> c1_n64_IO_out, 
            c1_n65_IO_out=> c1_n65_IO_out, 
            c1_n66_IO_out=> c1_n66_IO_out, 
            c1_n67_IO_out=> c1_n67_IO_out, 
            c1_n68_IO_out=> c1_n68_IO_out, 
            c1_n69_IO_out=> c1_n69_IO_out, 
            c1_n70_IO_out=> c1_n70_IO_out, 
            c1_n71_IO_out=> c1_n71_IO_out, 
            c1_n72_IO_out=> c1_n72_IO_out, 
            c1_n73_IO_out=> c1_n73_IO_out, 
            c1_n74_IO_out=> c1_n74_IO_out, 
            c1_n75_IO_out=> c1_n75_IO_out, 
            c1_n76_IO_out=> c1_n76_IO_out, 
            c1_n77_IO_out=> c1_n77_IO_out, 
            c1_n78_IO_out=> c1_n78_IO_out, 
            c1_n79_IO_out=> c1_n79_IO_out, 
            c1_n80_IO_out=> c1_n80_IO_out, 
            c1_n81_IO_out=> c1_n81_IO_out, 
            c1_n82_IO_out=> c1_n82_IO_out, 
            c1_n83_IO_out=> c1_n83_IO_out, 
            c1_n84_IO_out=> c1_n84_IO_out, 
            c1_n85_IO_out=> c1_n85_IO_out, 
            c1_n86_IO_out=> c1_n86_IO_out, 
            c1_n87_IO_out=> c1_n87_IO_out, 
            c1_n88_IO_out=> c1_n88_IO_out, 
            c1_n89_IO_out=> c1_n89_IO_out, 
            c1_n90_IO_out=> c1_n90_IO_out, 
            c1_n91_IO_out=> c1_n91_IO_out, 
            c1_n92_IO_out=> c1_n92_IO_out, 
            c1_n93_IO_out=> c1_n93_IO_out, 
            c1_n94_IO_out=> c1_n94_IO_out, 
            c1_n95_IO_out=> c1_n95_IO_out, 
            c1_n96_IO_out=> c1_n96_IO_out, 
            c1_n97_IO_out=> c1_n97_IO_out, 
            c1_n98_IO_out=> c1_n98_IO_out, 
            c1_n99_IO_out=> c1_n99_IO_out, 
            c1_n100_IO_out=> c1_n100_IO_out, 
            c1_n101_IO_out=> c1_n101_IO_out, 
            c1_n102_IO_out=> c1_n102_IO_out, 
            c1_n103_IO_out=> c1_n103_IO_out, 
            c1_n104_IO_out=> c1_n104_IO_out, 
            c1_n105_IO_out=> c1_n105_IO_out, 
            c1_n106_IO_out=> c1_n106_IO_out, 
            c1_n107_IO_out=> c1_n107_IO_out, 
            c1_n108_IO_out=> c1_n108_IO_out, 
            c1_n109_IO_out=> c1_n109_IO_out, 
            c1_n110_IO_out=> c1_n110_IO_out, 
            c1_n111_IO_out=> c1_n111_IO_out, 
            c1_n112_IO_out=> c1_n112_IO_out, 
            c1_n113_IO_out=> c1_n113_IO_out, 
            c1_n114_IO_out=> c1_n114_IO_out, 
            c1_n115_IO_out=> c1_n115_IO_out, 
            c1_n116_IO_out=> c1_n116_IO_out, 
            c1_n117_IO_out=> c1_n117_IO_out, 
            c1_n118_IO_out=> c1_n118_IO_out, 
            c1_n119_IO_out=> c1_n119_IO_out, 
            c1_n120_IO_out=> c1_n120_IO_out, 
            c1_n121_IO_out=> c1_n121_IO_out, 
            c1_n122_IO_out=> c1_n122_IO_out, 
            c1_n123_IO_out=> c1_n123_IO_out, 
            c1_n124_IO_out=> c1_n124_IO_out, 
            c1_n125_IO_out=> c1_n125_IO_out, 
            c1_n126_IO_out=> c1_n126_IO_out, 
            c1_n127_IO_out=> c1_n127_IO_out, 
            c1_n128_IO_out=> c1_n128_IO_out, 
            c1_n129_IO_out=> c1_n129_IO_out, 
            c1_n130_IO_out=> c1_n130_IO_out, 
            c1_n131_IO_out=> c1_n131_IO_out, 
            c1_n132_IO_out=> c1_n132_IO_out, 
            c1_n133_IO_out=> c1_n133_IO_out, 
            c1_n134_IO_out=> c1_n134_IO_out, 
            c1_n135_IO_out=> c1_n135_IO_out, 
            c1_n136_IO_out=> c1_n136_IO_out, 
            c1_n137_IO_out=> c1_n137_IO_out, 
            c1_n138_IO_out=> c1_n138_IO_out, 
            c1_n139_IO_out=> c1_n139_IO_out, 
            c1_n140_IO_out=> c1_n140_IO_out, 
            c1_n141_IO_out=> c1_n141_IO_out, 
            c1_n142_IO_out=> c1_n142_IO_out, 
            c1_n143_IO_out=> c1_n143_IO_out, 
            c1_n144_IO_out=> c1_n144_IO_out, 
            c1_n145_IO_out=> c1_n145_IO_out, 
            c1_n146_IO_out=> c1_n146_IO_out, 
            c1_n147_IO_out=> c1_n147_IO_out, 
            c1_n148_IO_out=> c1_n148_IO_out, 
            c1_n149_IO_out=> c1_n149_IO_out, 
            c1_n150_IO_out=> c1_n150_IO_out, 
            c1_n151_IO_out=> c1_n151_IO_out, 
            c1_n152_IO_out=> c1_n152_IO_out, 
            c1_n153_IO_out=> c1_n153_IO_out, 
            c1_n154_IO_out=> c1_n154_IO_out, 
            c1_n155_IO_out=> c1_n155_IO_out, 
            c1_n156_IO_out=> c1_n156_IO_out, 
            c1_n157_IO_out=> c1_n157_IO_out, 
            c1_n158_IO_out=> c1_n158_IO_out, 
            c1_n159_IO_out=> c1_n159_IO_out, 
            c1_n160_IO_out=> c1_n160_IO_out, 
            c1_n161_IO_out=> c1_n161_IO_out, 
            c1_n162_IO_out=> c1_n162_IO_out, 
            c1_n163_IO_out=> c1_n163_IO_out, 
            c1_n164_IO_out=> c1_n164_IO_out, 
            c1_n165_IO_out=> c1_n165_IO_out, 
            c1_n166_IO_out=> c1_n166_IO_out, 
            c1_n167_IO_out=> c1_n167_IO_out, 
            c1_n168_IO_out=> c1_n168_IO_out, 
            c1_n169_IO_out=> c1_n169_IO_out, 
            c1_n170_IO_out=> c1_n170_IO_out, 
            c1_n171_IO_out=> c1_n171_IO_out, 
            c1_n172_IO_out=> c1_n172_IO_out, 
            c1_n173_IO_out=> c1_n173_IO_out, 
            c1_n174_IO_out=> c1_n174_IO_out, 
            c1_n175_IO_out=> c1_n175_IO_out, 
            c1_n176_IO_out=> c1_n176_IO_out, 
            c1_n177_IO_out=> c1_n177_IO_out, 
            c1_n178_IO_out=> c1_n178_IO_out, 
            c1_n179_IO_out=> c1_n179_IO_out, 
            c1_n180_IO_out=> c1_n180_IO_out, 
            c1_n181_IO_out=> c1_n181_IO_out, 
            c1_n182_IO_out=> c1_n182_IO_out, 
            c1_n183_IO_out=> c1_n183_IO_out, 
            c1_n184_IO_out=> c1_n184_IO_out, 
            c1_n185_IO_out=> c1_n185_IO_out, 
            c1_n186_IO_out=> c1_n186_IO_out, 
            c1_n187_IO_out=> c1_n187_IO_out, 
            c1_n188_IO_out=> c1_n188_IO_out, 
            c1_n189_IO_out=> c1_n189_IO_out, 
            c1_n190_IO_out=> c1_n190_IO_out, 
            c1_n191_IO_out=> c1_n191_IO_out, 
            c1_n192_IO_out=> c1_n192_IO_out, 
            c1_n193_IO_out=> c1_n193_IO_out, 
            c1_n194_IO_out=> c1_n194_IO_out, 
            c1_n195_IO_out=> c1_n195_IO_out, 
            c1_n196_IO_out=> c1_n196_IO_out, 
            c1_n197_IO_out=> c1_n197_IO_out, 
            c1_n198_IO_out=> c1_n198_IO_out, 
            c1_n199_IO_out=> c1_n199_IO_out, 
            c1_n200_IO_out=> c1_n200_IO_out, 
            c1_n201_IO_out=> c1_n201_IO_out, 
            c1_n202_IO_out=> c1_n202_IO_out, 
            c1_n203_IO_out=> c1_n203_IO_out, 
            c1_n204_IO_out=> c1_n204_IO_out, 
            c1_n205_IO_out=> c1_n205_IO_out, 
            c1_n206_IO_out=> c1_n206_IO_out, 
            c1_n207_IO_out=> c1_n207_IO_out, 
            c1_n208_IO_out=> c1_n208_IO_out, 
            c1_n209_IO_out=> c1_n209_IO_out, 
            c1_n210_IO_out=> c1_n210_IO_out, 
            c1_n211_IO_out=> c1_n211_IO_out, 
            c1_n212_IO_out=> c1_n212_IO_out, 
            c1_n213_IO_out=> c1_n213_IO_out, 
            c1_n214_IO_out=> c1_n214_IO_out, 
            c1_n215_IO_out=> c1_n215_IO_out, 
            c1_n216_IO_out=> c1_n216_IO_out, 
            c1_n217_IO_out=> c1_n217_IO_out, 
            c1_n218_IO_out=> c1_n218_IO_out, 
            c1_n219_IO_out=> c1_n219_IO_out, 
            c1_n220_IO_out=> c1_n220_IO_out, 
            c1_n221_IO_out=> c1_n221_IO_out, 
            c1_n222_IO_out=> c1_n222_IO_out, 
            c1_n223_IO_out=> c1_n223_IO_out, 
            c1_n224_IO_out=> c1_n224_IO_out, 
            c1_n225_IO_out=> c1_n225_IO_out, 
            c1_n226_IO_out=> c1_n226_IO_out, 
            c1_n227_IO_out=> c1_n227_IO_out, 
            c1_n228_IO_out=> c1_n228_IO_out, 
            c1_n229_IO_out=> c1_n229_IO_out, 
            c1_n230_IO_out=> c1_n230_IO_out, 
            c1_n231_IO_out=> c1_n231_IO_out, 
            c1_n232_IO_out=> c1_n232_IO_out, 
            c1_n233_IO_out=> c1_n233_IO_out, 
            c1_n234_IO_out=> c1_n234_IO_out, 
            c1_n235_IO_out=> c1_n235_IO_out, 
            c1_n236_IO_out=> c1_n236_IO_out, 
            c1_n237_IO_out=> c1_n237_IO_out, 
            c1_n238_IO_out=> c1_n238_IO_out, 
            c1_n239_IO_out=> c1_n239_IO_out, 
            c1_n240_IO_out=> c1_n240_IO_out, 
            c1_n241_IO_out=> c1_n241_IO_out, 
            c1_n242_IO_out=> c1_n242_IO_out, 
            c1_n243_IO_out=> c1_n243_IO_out, 
            c1_n244_IO_out=> c1_n244_IO_out, 
            c1_n245_IO_out=> c1_n245_IO_out, 
            c1_n246_IO_out=> c1_n246_IO_out, 
            c1_n247_IO_out=> c1_n247_IO_out, 
            c1_n248_IO_out=> c1_n248_IO_out, 
            c1_n249_IO_out=> c1_n249_IO_out, 
            c1_n250_IO_out=> c1_n250_IO_out, 
            c1_n251_IO_out=> c1_n251_IO_out, 
            c1_n252_IO_out=> c1_n252_IO_out, 
            c1_n253_IO_out=> c1_n253_IO_out, 
            c1_n254_IO_out=> c1_n254_IO_out, 
            c1_n255_IO_out=> c1_n255_IO_out, 
            c1_n256_IO_out=> c1_n256_IO_out, 
            c1_n257_IO_out=> c1_n257_IO_out, 
            c1_n258_IO_out=> c1_n258_IO_out, 
            c1_n259_IO_out=> c1_n259_IO_out, 
            c1_n260_IO_out=> c1_n260_IO_out, 
            c1_n261_IO_out=> c1_n261_IO_out, 
            c1_n262_IO_out=> c1_n262_IO_out, 
            c1_n263_IO_out=> c1_n263_IO_out, 
            c1_n264_IO_out=> c1_n264_IO_out, 
            c1_n265_IO_out=> c1_n265_IO_out, 
            c1_n266_IO_out=> c1_n266_IO_out, 
            c1_n267_IO_out=> c1_n267_IO_out, 
            c1_n268_IO_out=> c1_n268_IO_out, 
            c1_n269_IO_out=> c1_n269_IO_out, 
            c1_n270_IO_out=> c1_n270_IO_out, 
            c1_n271_IO_out=> c1_n271_IO_out, 
            c1_n272_IO_out=> c1_n272_IO_out, 
            c1_n273_IO_out=> c1_n273_IO_out, 
            c1_n274_IO_out=> c1_n274_IO_out, 
            c1_n275_IO_out=> c1_n275_IO_out, 
            c1_n276_IO_out=> c1_n276_IO_out, 
            c1_n277_IO_out=> c1_n277_IO_out, 
            c1_n278_IO_out=> c1_n278_IO_out, 
            c1_n279_IO_out=> c1_n279_IO_out, 
            c1_n280_IO_out=> c1_n280_IO_out, 
            c1_n281_IO_out=> c1_n281_IO_out, 
            c1_n282_IO_out=> c1_n282_IO_out, 
            c1_n283_IO_out=> c1_n283_IO_out, 
            c1_n284_IO_out=> c1_n284_IO_out, 
            c1_n285_IO_out=> c1_n285_IO_out, 
            c1_n286_IO_out=> c1_n286_IO_out, 
            c1_n287_IO_out=> c1_n287_IO_out, 
            c1_n288_IO_out=> c1_n288_IO_out, 
            c1_n289_IO_out=> c1_n289_IO_out, 
            c1_n290_IO_out=> c1_n290_IO_out, 
            c1_n291_IO_out=> c1_n291_IO_out, 
            c1_n292_IO_out=> c1_n292_IO_out, 
            c1_n293_IO_out=> c1_n293_IO_out, 
            c1_n294_IO_out=> c1_n294_IO_out, 
            c1_n295_IO_out=> c1_n295_IO_out, 
            c1_n296_IO_out=> c1_n296_IO_out, 
            c1_n297_IO_out=> c1_n297_IO_out, 
            c1_n298_IO_out=> c1_n298_IO_out, 
            c1_n299_IO_out=> c1_n299_IO_out, 
            -- ['OUT']['manual'] 
            c1_n0_W_out=> c1_n0_W_out, 
            c1_n1_W_out=> c1_n1_W_out, 
            c1_n2_W_out=> c1_n2_W_out, 
            c1_n3_W_out=> c1_n3_W_out, 
            c1_n4_W_out=> c1_n4_W_out, 
            c1_n5_W_out=> c1_n5_W_out, 
            c1_n6_W_out=> c1_n6_W_out, 
            c1_n7_W_out=> c1_n7_W_out, 
            c1_n8_W_out=> c1_n8_W_out, 
            c1_n9_W_out=> c1_n9_W_out, 
            c1_n10_W_out=> c1_n10_W_out, 
            c1_n11_W_out=> c1_n11_W_out, 
            c1_n12_W_out=> c1_n12_W_out, 
            c1_n13_W_out=> c1_n13_W_out, 
            c1_n14_W_out=> c1_n14_W_out, 
            c1_n15_W_out=> c1_n15_W_out, 
            c1_n16_W_out=> c1_n16_W_out, 
            c1_n17_W_out=> c1_n17_W_out, 
            c1_n18_W_out=> c1_n18_W_out, 
            c1_n19_W_out=> c1_n19_W_out, 
            c1_n20_W_out=> c1_n20_W_out, 
            c1_n21_W_out=> c1_n21_W_out, 
            c1_n22_W_out=> c1_n22_W_out, 
            c1_n23_W_out=> c1_n23_W_out, 
            c1_n24_W_out=> c1_n24_W_out, 
            c1_n25_W_out=> c1_n25_W_out, 
            c1_n26_W_out=> c1_n26_W_out, 
            c1_n27_W_out=> c1_n27_W_out, 
            c1_n28_W_out=> c1_n28_W_out, 
            c1_n29_W_out=> c1_n29_W_out, 
            c1_n30_W_out=> c1_n30_W_out, 
            c1_n31_W_out=> c1_n31_W_out, 
            c1_n32_W_out=> c1_n32_W_out, 
            c1_n33_W_out=> c1_n33_W_out, 
            c1_n34_W_out=> c1_n34_W_out, 
            c1_n35_W_out=> c1_n35_W_out, 
            c1_n36_W_out=> c1_n36_W_out, 
            c1_n37_W_out=> c1_n37_W_out, 
            c1_n38_W_out=> c1_n38_W_out, 
            c1_n39_W_out=> c1_n39_W_out, 
            c1_n40_W_out=> c1_n40_W_out, 
            c1_n41_W_out=> c1_n41_W_out, 
            c1_n42_W_out=> c1_n42_W_out, 
            c1_n43_W_out=> c1_n43_W_out, 
            c1_n44_W_out=> c1_n44_W_out, 
            c1_n45_W_out=> c1_n45_W_out, 
            c1_n46_W_out=> c1_n46_W_out, 
            c1_n47_W_out=> c1_n47_W_out, 
            c1_n48_W_out=> c1_n48_W_out, 
            c1_n49_W_out=> c1_n49_W_out, 
            c1_n50_W_out=> c1_n50_W_out, 
            c1_n51_W_out=> c1_n51_W_out, 
            c1_n52_W_out=> c1_n52_W_out, 
            c1_n53_W_out=> c1_n53_W_out, 
            c1_n54_W_out=> c1_n54_W_out, 
            c1_n55_W_out=> c1_n55_W_out, 
            c1_n56_W_out=> c1_n56_W_out, 
            c1_n57_W_out=> c1_n57_W_out, 
            c1_n58_W_out=> c1_n58_W_out, 
            c1_n59_W_out=> c1_n59_W_out, 
            c1_n60_W_out=> c1_n60_W_out, 
            c1_n61_W_out=> c1_n61_W_out, 
            c1_n62_W_out=> c1_n62_W_out, 
            c1_n63_W_out=> c1_n63_W_out, 
            c1_n64_W_out=> c1_n64_W_out, 
            c1_n65_W_out=> c1_n65_W_out, 
            c1_n66_W_out=> c1_n66_W_out, 
            c1_n67_W_out=> c1_n67_W_out, 
            c1_n68_W_out=> c1_n68_W_out, 
            c1_n69_W_out=> c1_n69_W_out, 
            c1_n70_W_out=> c1_n70_W_out, 
            c1_n71_W_out=> c1_n71_W_out, 
            c1_n72_W_out=> c1_n72_W_out, 
            c1_n73_W_out=> c1_n73_W_out, 
            c1_n74_W_out=> c1_n74_W_out, 
            c1_n75_W_out=> c1_n75_W_out, 
            c1_n76_W_out=> c1_n76_W_out, 
            c1_n77_W_out=> c1_n77_W_out, 
            c1_n78_W_out=> c1_n78_W_out, 
            c1_n79_W_out=> c1_n79_W_out, 
            c1_n80_W_out=> c1_n80_W_out, 
            c1_n81_W_out=> c1_n81_W_out, 
            c1_n82_W_out=> c1_n82_W_out, 
            c1_n83_W_out=> c1_n83_W_out, 
            c1_n84_W_out=> c1_n84_W_out, 
            c1_n85_W_out=> c1_n85_W_out, 
            c1_n86_W_out=> c1_n86_W_out, 
            c1_n87_W_out=> c1_n87_W_out, 
            c1_n88_W_out=> c1_n88_W_out, 
            c1_n89_W_out=> c1_n89_W_out, 
            c1_n90_W_out=> c1_n90_W_out, 
            c1_n91_W_out=> c1_n91_W_out, 
            c1_n92_W_out=> c1_n92_W_out, 
            c1_n93_W_out=> c1_n93_W_out, 
            c1_n94_W_out=> c1_n94_W_out, 
            c1_n95_W_out=> c1_n95_W_out, 
            c1_n96_W_out=> c1_n96_W_out, 
            c1_n97_W_out=> c1_n97_W_out, 
            c1_n98_W_out=> c1_n98_W_out, 
            c1_n99_W_out=> c1_n99_W_out, 
            c1_n100_W_out=> c1_n100_W_out, 
            c1_n101_W_out=> c1_n101_W_out, 
            c1_n102_W_out=> c1_n102_W_out, 
            c1_n103_W_out=> c1_n103_W_out, 
            c1_n104_W_out=> c1_n104_W_out, 
            c1_n105_W_out=> c1_n105_W_out, 
            c1_n106_W_out=> c1_n106_W_out, 
            c1_n107_W_out=> c1_n107_W_out, 
            c1_n108_W_out=> c1_n108_W_out, 
            c1_n109_W_out=> c1_n109_W_out, 
            c1_n110_W_out=> c1_n110_W_out, 
            c1_n111_W_out=> c1_n111_W_out, 
            c1_n112_W_out=> c1_n112_W_out, 
            c1_n113_W_out=> c1_n113_W_out, 
            c1_n114_W_out=> c1_n114_W_out, 
            c1_n115_W_out=> c1_n115_W_out, 
            c1_n116_W_out=> c1_n116_W_out, 
            c1_n117_W_out=> c1_n117_W_out, 
            c1_n118_W_out=> c1_n118_W_out, 
            c1_n119_W_out=> c1_n119_W_out, 
            c1_n120_W_out=> c1_n120_W_out, 
            c1_n121_W_out=> c1_n121_W_out, 
            c1_n122_W_out=> c1_n122_W_out, 
            c1_n123_W_out=> c1_n123_W_out, 
            c1_n124_W_out=> c1_n124_W_out, 
            c1_n125_W_out=> c1_n125_W_out, 
            c1_n126_W_out=> c1_n126_W_out, 
            c1_n127_W_out=> c1_n127_W_out, 
            c1_n128_W_out=> c1_n128_W_out, 
            c1_n129_W_out=> c1_n129_W_out, 
            c1_n130_W_out=> c1_n130_W_out, 
            c1_n131_W_out=> c1_n131_W_out, 
            c1_n132_W_out=> c1_n132_W_out, 
            c1_n133_W_out=> c1_n133_W_out, 
            c1_n134_W_out=> c1_n134_W_out, 
            c1_n135_W_out=> c1_n135_W_out, 
            c1_n136_W_out=> c1_n136_W_out, 
            c1_n137_W_out=> c1_n137_W_out, 
            c1_n138_W_out=> c1_n138_W_out, 
            c1_n139_W_out=> c1_n139_W_out, 
            c1_n140_W_out=> c1_n140_W_out, 
            c1_n141_W_out=> c1_n141_W_out, 
            c1_n142_W_out=> c1_n142_W_out, 
            c1_n143_W_out=> c1_n143_W_out, 
            c1_n144_W_out=> c1_n144_W_out, 
            c1_n145_W_out=> c1_n145_W_out, 
            c1_n146_W_out=> c1_n146_W_out, 
            c1_n147_W_out=> c1_n147_W_out, 
            c1_n148_W_out=> c1_n148_W_out, 
            c1_n149_W_out=> c1_n149_W_out, 
            c1_n150_W_out=> c1_n150_W_out, 
            c1_n151_W_out=> c1_n151_W_out, 
            c1_n152_W_out=> c1_n152_W_out, 
            c1_n153_W_out=> c1_n153_W_out, 
            c1_n154_W_out=> c1_n154_W_out, 
            c1_n155_W_out=> c1_n155_W_out, 
            c1_n156_W_out=> c1_n156_W_out, 
            c1_n157_W_out=> c1_n157_W_out, 
            c1_n158_W_out=> c1_n158_W_out, 
            c1_n159_W_out=> c1_n159_W_out, 
            c1_n160_W_out=> c1_n160_W_out, 
            c1_n161_W_out=> c1_n161_W_out, 
            c1_n162_W_out=> c1_n162_W_out, 
            c1_n163_W_out=> c1_n163_W_out, 
            c1_n164_W_out=> c1_n164_W_out, 
            c1_n165_W_out=> c1_n165_W_out, 
            c1_n166_W_out=> c1_n166_W_out, 
            c1_n167_W_out=> c1_n167_W_out, 
            c1_n168_W_out=> c1_n168_W_out, 
            c1_n169_W_out=> c1_n169_W_out, 
            c1_n170_W_out=> c1_n170_W_out, 
            c1_n171_W_out=> c1_n171_W_out, 
            c1_n172_W_out=> c1_n172_W_out, 
            c1_n173_W_out=> c1_n173_W_out, 
            c1_n174_W_out=> c1_n174_W_out, 
            c1_n175_W_out=> c1_n175_W_out, 
            c1_n176_W_out=> c1_n176_W_out, 
            c1_n177_W_out=> c1_n177_W_out, 
            c1_n178_W_out=> c1_n178_W_out, 
            c1_n179_W_out=> c1_n179_W_out, 
            c1_n180_W_out=> c1_n180_W_out, 
            c1_n181_W_out=> c1_n181_W_out, 
            c1_n182_W_out=> c1_n182_W_out, 
            c1_n183_W_out=> c1_n183_W_out, 
            c1_n184_W_out=> c1_n184_W_out, 
            c1_n185_W_out=> c1_n185_W_out, 
            c1_n186_W_out=> c1_n186_W_out, 
            c1_n187_W_out=> c1_n187_W_out, 
            c1_n188_W_out=> c1_n188_W_out, 
            c1_n189_W_out=> c1_n189_W_out, 
            c1_n190_W_out=> c1_n190_W_out, 
            c1_n191_W_out=> c1_n191_W_out, 
            c1_n192_W_out=> c1_n192_W_out, 
            c1_n193_W_out=> c1_n193_W_out, 
            c1_n194_W_out=> c1_n194_W_out, 
            c1_n195_W_out=> c1_n195_W_out, 
            c1_n196_W_out=> c1_n196_W_out, 
            c1_n197_W_out=> c1_n197_W_out, 
            c1_n198_W_out=> c1_n198_W_out, 
            c1_n199_W_out=> c1_n199_W_out, 
            c1_n200_W_out=> c1_n200_W_out, 
            c1_n201_W_out=> c1_n201_W_out, 
            c1_n202_W_out=> c1_n202_W_out, 
            c1_n203_W_out=> c1_n203_W_out, 
            c1_n204_W_out=> c1_n204_W_out, 
            c1_n205_W_out=> c1_n205_W_out, 
            c1_n206_W_out=> c1_n206_W_out, 
            c1_n207_W_out=> c1_n207_W_out, 
            c1_n208_W_out=> c1_n208_W_out, 
            c1_n209_W_out=> c1_n209_W_out, 
            c1_n210_W_out=> c1_n210_W_out, 
            c1_n211_W_out=> c1_n211_W_out, 
            c1_n212_W_out=> c1_n212_W_out, 
            c1_n213_W_out=> c1_n213_W_out, 
            c1_n214_W_out=> c1_n214_W_out, 
            c1_n215_W_out=> c1_n215_W_out, 
            c1_n216_W_out=> c1_n216_W_out, 
            c1_n217_W_out=> c1_n217_W_out, 
            c1_n218_W_out=> c1_n218_W_out, 
            c1_n219_W_out=> c1_n219_W_out, 
            c1_n220_W_out=> c1_n220_W_out, 
            c1_n221_W_out=> c1_n221_W_out, 
            c1_n222_W_out=> c1_n222_W_out, 
            c1_n223_W_out=> c1_n223_W_out, 
            c1_n224_W_out=> c1_n224_W_out, 
            c1_n225_W_out=> c1_n225_W_out, 
            c1_n226_W_out=> c1_n226_W_out, 
            c1_n227_W_out=> c1_n227_W_out, 
            c1_n228_W_out=> c1_n228_W_out, 
            c1_n229_W_out=> c1_n229_W_out, 
            c1_n230_W_out=> c1_n230_W_out, 
            c1_n231_W_out=> c1_n231_W_out, 
            c1_n232_W_out=> c1_n232_W_out, 
            c1_n233_W_out=> c1_n233_W_out, 
            c1_n234_W_out=> c1_n234_W_out, 
            c1_n235_W_out=> c1_n235_W_out, 
            c1_n236_W_out=> c1_n236_W_out, 
            c1_n237_W_out=> c1_n237_W_out, 
            c1_n238_W_out=> c1_n238_W_out, 
            c1_n239_W_out=> c1_n239_W_out, 
            c1_n240_W_out=> c1_n240_W_out, 
            c1_n241_W_out=> c1_n241_W_out, 
            c1_n242_W_out=> c1_n242_W_out, 
            c1_n243_W_out=> c1_n243_W_out, 
            c1_n244_W_out=> c1_n244_W_out, 
            c1_n245_W_out=> c1_n245_W_out, 
            c1_n246_W_out=> c1_n246_W_out, 
            c1_n247_W_out=> c1_n247_W_out, 
            c1_n248_W_out=> c1_n248_W_out, 
            c1_n249_W_out=> c1_n249_W_out, 
            c1_n250_W_out=> c1_n250_W_out, 
            c1_n251_W_out=> c1_n251_W_out, 
            c1_n252_W_out=> c1_n252_W_out, 
            c1_n253_W_out=> c1_n253_W_out, 
            c1_n254_W_out=> c1_n254_W_out, 
            c1_n255_W_out=> c1_n255_W_out, 
            c1_n256_W_out=> c1_n256_W_out, 
            c1_n257_W_out=> c1_n257_W_out, 
            c1_n258_W_out=> c1_n258_W_out, 
            c1_n259_W_out=> c1_n259_W_out, 
            c1_n260_W_out=> c1_n260_W_out, 
            c1_n261_W_out=> c1_n261_W_out, 
            c1_n262_W_out=> c1_n262_W_out, 
            c1_n263_W_out=> c1_n263_W_out, 
            c1_n264_W_out=> c1_n264_W_out, 
            c1_n265_W_out=> c1_n265_W_out, 
            c1_n266_W_out=> c1_n266_W_out, 
            c1_n267_W_out=> c1_n267_W_out, 
            c1_n268_W_out=> c1_n268_W_out, 
            c1_n269_W_out=> c1_n269_W_out, 
            c1_n270_W_out=> c1_n270_W_out, 
            c1_n271_W_out=> c1_n271_W_out, 
            c1_n272_W_out=> c1_n272_W_out, 
            c1_n273_W_out=> c1_n273_W_out, 
            c1_n274_W_out=> c1_n274_W_out, 
            c1_n275_W_out=> c1_n275_W_out, 
            c1_n276_W_out=> c1_n276_W_out, 
            c1_n277_W_out=> c1_n277_W_out, 
            c1_n278_W_out=> c1_n278_W_out, 
            c1_n279_W_out=> c1_n279_W_out, 
            c1_n280_W_out=> c1_n280_W_out, 
            c1_n281_W_out=> c1_n281_W_out, 
            c1_n282_W_out=> c1_n282_W_out, 
            c1_n283_W_out=> c1_n283_W_out, 
            c1_n284_W_out=> c1_n284_W_out, 
            c1_n285_W_out=> c1_n285_W_out, 
            c1_n286_W_out=> c1_n286_W_out, 
            c1_n287_W_out=> c1_n287_W_out, 
            c1_n288_W_out=> c1_n288_W_out, 
            c1_n289_W_out=> c1_n289_W_out, 
            c1_n290_W_out=> c1_n290_W_out, 
            c1_n291_W_out=> c1_n291_W_out, 
            c1_n292_W_out=> c1_n292_W_out, 
            c1_n293_W_out=> c1_n293_W_out, 
            c1_n294_W_out=> c1_n294_W_out, 
            c1_n295_W_out=> c1_n295_W_out, 
            c1_n296_W_out=> c1_n296_W_out, 
            c1_n297_W_out=> c1_n297_W_out, 
            c1_n298_W_out=> c1_n298_W_out, 
            c1_n299_W_out=> c1_n299_W_out
   );
            
camada2_inst_2: ENTITY work.camada2_ReLU_100neuron_8bits_300n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c2_IO_in, 
            c2_n0_W_in=> c1_n0_W_out,
            c2_n1_W_in=> c1_n1_W_out,
            c2_n2_W_in=> c1_n2_W_out,
            c2_n3_W_in=> c1_n3_W_out,
            c2_n4_W_in=> c1_n4_W_out,
            c2_n5_W_in=> c1_n5_W_out,
            c2_n6_W_in=> c1_n6_W_out,
            c2_n7_W_in=> c1_n7_W_out,
            c2_n8_W_in=> c1_n8_W_out,
            c2_n9_W_in=> c1_n9_W_out,
            c2_n10_W_in=> c1_n10_W_out,
            c2_n11_W_in=> c1_n11_W_out,
            c2_n12_W_in=> c1_n12_W_out,
            c2_n13_W_in=> c1_n13_W_out,
            c2_n14_W_in=> c1_n14_W_out,
            c2_n15_W_in=> c1_n15_W_out,
            c2_n16_W_in=> c1_n16_W_out,
            c2_n17_W_in=> c1_n17_W_out,
            c2_n18_W_in=> c1_n18_W_out,
            c2_n19_W_in=> c1_n19_W_out,
            c2_n20_W_in=> c1_n20_W_out,
            c2_n21_W_in=> c1_n21_W_out,
            c2_n22_W_in=> c1_n22_W_out,
            c2_n23_W_in=> c1_n23_W_out,
            c2_n24_W_in=> c1_n24_W_out,
            c2_n25_W_in=> c1_n25_W_out,
            c2_n26_W_in=> c1_n26_W_out,
            c2_n27_W_in=> c1_n27_W_out,
            c2_n28_W_in=> c1_n28_W_out,
            c2_n29_W_in=> c1_n29_W_out,
            c2_n30_W_in=> c1_n30_W_out,
            c2_n31_W_in=> c1_n31_W_out,
            c2_n32_W_in=> c1_n32_W_out,
            c2_n33_W_in=> c1_n33_W_out,
            c2_n34_W_in=> c1_n34_W_out,
            c2_n35_W_in=> c1_n35_W_out,
            c2_n36_W_in=> c1_n36_W_out,
            c2_n37_W_in=> c1_n37_W_out,
            c2_n38_W_in=> c1_n38_W_out,
            c2_n39_W_in=> c1_n39_W_out,
            c2_n40_W_in=> c1_n40_W_out,
            c2_n41_W_in=> c1_n41_W_out,
            c2_n42_W_in=> c1_n42_W_out,
            c2_n43_W_in=> c1_n43_W_out,
            c2_n44_W_in=> c1_n44_W_out,
            c2_n45_W_in=> c1_n45_W_out,
            c2_n46_W_in=> c1_n46_W_out,
            c2_n47_W_in=> c1_n47_W_out,
            c2_n48_W_in=> c1_n48_W_out,
            c2_n49_W_in=> c1_n49_W_out,
            c2_n50_W_in=> c1_n50_W_out,
            c2_n51_W_in=> c1_n51_W_out,
            c2_n52_W_in=> c1_n52_W_out,
            c2_n53_W_in=> c1_n53_W_out,
            c2_n54_W_in=> c1_n54_W_out,
            c2_n55_W_in=> c1_n55_W_out,
            c2_n56_W_in=> c1_n56_W_out,
            c2_n57_W_in=> c1_n57_W_out,
            c2_n58_W_in=> c1_n58_W_out,
            c2_n59_W_in=> c1_n59_W_out,
            c2_n60_W_in=> c1_n60_W_out,
            c2_n61_W_in=> c1_n61_W_out,
            c2_n62_W_in=> c1_n62_W_out,
            c2_n63_W_in=> c1_n63_W_out,
            c2_n64_W_in=> c1_n64_W_out,
            c2_n65_W_in=> c1_n65_W_out,
            c2_n66_W_in=> c1_n66_W_out,
            c2_n67_W_in=> c1_n67_W_out,
            c2_n68_W_in=> c1_n68_W_out,
            c2_n69_W_in=> c1_n69_W_out,
            c2_n70_W_in=> c1_n70_W_out,
            c2_n71_W_in=> c1_n71_W_out,
            c2_n72_W_in=> c1_n72_W_out,
            c2_n73_W_in=> c1_n73_W_out,
            c2_n74_W_in=> c1_n74_W_out,
            c2_n75_W_in=> c1_n75_W_out,
            c2_n76_W_in=> c1_n76_W_out,
            c2_n77_W_in=> c1_n77_W_out,
            c2_n78_W_in=> c1_n78_W_out,
            c2_n79_W_in=> c1_n79_W_out,
            c2_n80_W_in=> c1_n80_W_out,
            c2_n81_W_in=> c1_n81_W_out,
            c2_n82_W_in=> c1_n82_W_out,
            c2_n83_W_in=> c1_n83_W_out,
            c2_n84_W_in=> c1_n84_W_out,
            c2_n85_W_in=> c1_n85_W_out,
            c2_n86_W_in=> c1_n86_W_out,
            c2_n87_W_in=> c1_n87_W_out,
            c2_n88_W_in=> c1_n88_W_out,
            c2_n89_W_in=> c1_n89_W_out,
            c2_n90_W_in=> c1_n90_W_out,
            c2_n91_W_in=> c1_n91_W_out,
            c2_n92_W_in=> c1_n92_W_out,
            c2_n93_W_in=> c1_n93_W_out,
            c2_n94_W_in=> c1_n94_W_out,
            c2_n95_W_in=> c1_n95_W_out,
            c2_n96_W_in=> c1_n96_W_out,
            c2_n97_W_in=> c1_n97_W_out,
            c2_n98_W_in=> c1_n98_W_out,
            c2_n99_W_in=> c1_n99_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c2_n0_IO_out=> c2_n0_IO_out, 
            c2_n1_IO_out=> c2_n1_IO_out, 
            c2_n2_IO_out=> c2_n2_IO_out, 
            c2_n3_IO_out=> c2_n3_IO_out, 
            c2_n4_IO_out=> c2_n4_IO_out, 
            c2_n5_IO_out=> c2_n5_IO_out, 
            c2_n6_IO_out=> c2_n6_IO_out, 
            c2_n7_IO_out=> c2_n7_IO_out, 
            c2_n8_IO_out=> c2_n8_IO_out, 
            c2_n9_IO_out=> c2_n9_IO_out, 
            c2_n10_IO_out=> c2_n10_IO_out, 
            c2_n11_IO_out=> c2_n11_IO_out, 
            c2_n12_IO_out=> c2_n12_IO_out, 
            c2_n13_IO_out=> c2_n13_IO_out, 
            c2_n14_IO_out=> c2_n14_IO_out, 
            c2_n15_IO_out=> c2_n15_IO_out, 
            c2_n16_IO_out=> c2_n16_IO_out, 
            c2_n17_IO_out=> c2_n17_IO_out, 
            c2_n18_IO_out=> c2_n18_IO_out, 
            c2_n19_IO_out=> c2_n19_IO_out, 
            c2_n20_IO_out=> c2_n20_IO_out, 
            c2_n21_IO_out=> c2_n21_IO_out, 
            c2_n22_IO_out=> c2_n22_IO_out, 
            c2_n23_IO_out=> c2_n23_IO_out, 
            c2_n24_IO_out=> c2_n24_IO_out, 
            c2_n25_IO_out=> c2_n25_IO_out, 
            c2_n26_IO_out=> c2_n26_IO_out, 
            c2_n27_IO_out=> c2_n27_IO_out, 
            c2_n28_IO_out=> c2_n28_IO_out, 
            c2_n29_IO_out=> c2_n29_IO_out, 
            c2_n30_IO_out=> c2_n30_IO_out, 
            c2_n31_IO_out=> c2_n31_IO_out, 
            c2_n32_IO_out=> c2_n32_IO_out, 
            c2_n33_IO_out=> c2_n33_IO_out, 
            c2_n34_IO_out=> c2_n34_IO_out, 
            c2_n35_IO_out=> c2_n35_IO_out, 
            c2_n36_IO_out=> c2_n36_IO_out, 
            c2_n37_IO_out=> c2_n37_IO_out, 
            c2_n38_IO_out=> c2_n38_IO_out, 
            c2_n39_IO_out=> c2_n39_IO_out, 
            c2_n40_IO_out=> c2_n40_IO_out, 
            c2_n41_IO_out=> c2_n41_IO_out, 
            c2_n42_IO_out=> c2_n42_IO_out, 
            c2_n43_IO_out=> c2_n43_IO_out, 
            c2_n44_IO_out=> c2_n44_IO_out, 
            c2_n45_IO_out=> c2_n45_IO_out, 
            c2_n46_IO_out=> c2_n46_IO_out, 
            c2_n47_IO_out=> c2_n47_IO_out, 
            c2_n48_IO_out=> c2_n48_IO_out, 
            c2_n49_IO_out=> c2_n49_IO_out, 
            c2_n50_IO_out=> c2_n50_IO_out, 
            c2_n51_IO_out=> c2_n51_IO_out, 
            c2_n52_IO_out=> c2_n52_IO_out, 
            c2_n53_IO_out=> c2_n53_IO_out, 
            c2_n54_IO_out=> c2_n54_IO_out, 
            c2_n55_IO_out=> c2_n55_IO_out, 
            c2_n56_IO_out=> c2_n56_IO_out, 
            c2_n57_IO_out=> c2_n57_IO_out, 
            c2_n58_IO_out=> c2_n58_IO_out, 
            c2_n59_IO_out=> c2_n59_IO_out, 
            c2_n60_IO_out=> c2_n60_IO_out, 
            c2_n61_IO_out=> c2_n61_IO_out, 
            c2_n62_IO_out=> c2_n62_IO_out, 
            c2_n63_IO_out=> c2_n63_IO_out, 
            c2_n64_IO_out=> c2_n64_IO_out, 
            c2_n65_IO_out=> c2_n65_IO_out, 
            c2_n66_IO_out=> c2_n66_IO_out, 
            c2_n67_IO_out=> c2_n67_IO_out, 
            c2_n68_IO_out=> c2_n68_IO_out, 
            c2_n69_IO_out=> c2_n69_IO_out, 
            c2_n70_IO_out=> c2_n70_IO_out, 
            c2_n71_IO_out=> c2_n71_IO_out, 
            c2_n72_IO_out=> c2_n72_IO_out, 
            c2_n73_IO_out=> c2_n73_IO_out, 
            c2_n74_IO_out=> c2_n74_IO_out, 
            c2_n75_IO_out=> c2_n75_IO_out, 
            c2_n76_IO_out=> c2_n76_IO_out, 
            c2_n77_IO_out=> c2_n77_IO_out, 
            c2_n78_IO_out=> c2_n78_IO_out, 
            c2_n79_IO_out=> c2_n79_IO_out, 
            c2_n80_IO_out=> c2_n80_IO_out, 
            c2_n81_IO_out=> c2_n81_IO_out, 
            c2_n82_IO_out=> c2_n82_IO_out, 
            c2_n83_IO_out=> c2_n83_IO_out, 
            c2_n84_IO_out=> c2_n84_IO_out, 
            c2_n85_IO_out=> c2_n85_IO_out, 
            c2_n86_IO_out=> c2_n86_IO_out, 
            c2_n87_IO_out=> c2_n87_IO_out, 
            c2_n88_IO_out=> c2_n88_IO_out, 
            c2_n89_IO_out=> c2_n89_IO_out, 
            c2_n90_IO_out=> c2_n90_IO_out, 
            c2_n91_IO_out=> c2_n91_IO_out, 
            c2_n92_IO_out=> c2_n92_IO_out, 
            c2_n93_IO_out=> c2_n93_IO_out, 
            c2_n94_IO_out=> c2_n94_IO_out, 
            c2_n95_IO_out=> c2_n95_IO_out, 
            c2_n96_IO_out=> c2_n96_IO_out, 
            c2_n97_IO_out=> c2_n97_IO_out, 
            c2_n98_IO_out=> c2_n98_IO_out, 
            c2_n99_IO_out=> c2_n99_IO_out, 
            -- ['OUT']['manual'] 
            c2_n0_W_out=> c2_n0_W_out, 
            c2_n1_W_out=> c2_n1_W_out, 
            c2_n2_W_out=> c2_n2_W_out, 
            c2_n3_W_out=> c2_n3_W_out, 
            c2_n4_W_out=> c2_n4_W_out, 
            c2_n5_W_out=> c2_n5_W_out, 
            c2_n6_W_out=> c2_n6_W_out, 
            c2_n7_W_out=> c2_n7_W_out, 
            c2_n8_W_out=> c2_n8_W_out, 
            c2_n9_W_out=> c2_n9_W_out, 
            c2_n10_W_out=> c2_n10_W_out, 
            c2_n11_W_out=> c2_n11_W_out, 
            c2_n12_W_out=> c2_n12_W_out, 
            c2_n13_W_out=> c2_n13_W_out, 
            c2_n14_W_out=> c2_n14_W_out, 
            c2_n15_W_out=> c2_n15_W_out, 
            c2_n16_W_out=> c2_n16_W_out, 
            c2_n17_W_out=> c2_n17_W_out, 
            c2_n18_W_out=> c2_n18_W_out, 
            c2_n19_W_out=> c2_n19_W_out, 
            c2_n20_W_out=> c2_n20_W_out, 
            c2_n21_W_out=> c2_n21_W_out, 
            c2_n22_W_out=> c2_n22_W_out, 
            c2_n23_W_out=> c2_n23_W_out, 
            c2_n24_W_out=> c2_n24_W_out, 
            c2_n25_W_out=> c2_n25_W_out, 
            c2_n26_W_out=> c2_n26_W_out, 
            c2_n27_W_out=> c2_n27_W_out, 
            c2_n28_W_out=> c2_n28_W_out, 
            c2_n29_W_out=> c2_n29_W_out, 
            c2_n30_W_out=> c2_n30_W_out, 
            c2_n31_W_out=> c2_n31_W_out, 
            c2_n32_W_out=> c2_n32_W_out, 
            c2_n33_W_out=> c2_n33_W_out, 
            c2_n34_W_out=> c2_n34_W_out, 
            c2_n35_W_out=> c2_n35_W_out, 
            c2_n36_W_out=> c2_n36_W_out, 
            c2_n37_W_out=> c2_n37_W_out, 
            c2_n38_W_out=> c2_n38_W_out, 
            c2_n39_W_out=> c2_n39_W_out, 
            c2_n40_W_out=> c2_n40_W_out, 
            c2_n41_W_out=> c2_n41_W_out, 
            c2_n42_W_out=> c2_n42_W_out, 
            c2_n43_W_out=> c2_n43_W_out, 
            c2_n44_W_out=> c2_n44_W_out, 
            c2_n45_W_out=> c2_n45_W_out, 
            c2_n46_W_out=> c2_n46_W_out, 
            c2_n47_W_out=> c2_n47_W_out, 
            c2_n48_W_out=> c2_n48_W_out, 
            c2_n49_W_out=> c2_n49_W_out, 
            c2_n50_W_out=> c2_n50_W_out, 
            c2_n51_W_out=> c2_n51_W_out, 
            c2_n52_W_out=> c2_n52_W_out, 
            c2_n53_W_out=> c2_n53_W_out, 
            c2_n54_W_out=> c2_n54_W_out, 
            c2_n55_W_out=> c2_n55_W_out, 
            c2_n56_W_out=> c2_n56_W_out, 
            c2_n57_W_out=> c2_n57_W_out, 
            c2_n58_W_out=> c2_n58_W_out, 
            c2_n59_W_out=> c2_n59_W_out, 
            c2_n60_W_out=> c2_n60_W_out, 
            c2_n61_W_out=> c2_n61_W_out, 
            c2_n62_W_out=> c2_n62_W_out, 
            c2_n63_W_out=> c2_n63_W_out, 
            c2_n64_W_out=> c2_n64_W_out, 
            c2_n65_W_out=> c2_n65_W_out, 
            c2_n66_W_out=> c2_n66_W_out, 
            c2_n67_W_out=> c2_n67_W_out, 
            c2_n68_W_out=> c2_n68_W_out, 
            c2_n69_W_out=> c2_n69_W_out, 
            c2_n70_W_out=> c2_n70_W_out, 
            c2_n71_W_out=> c2_n71_W_out, 
            c2_n72_W_out=> c2_n72_W_out, 
            c2_n73_W_out=> c2_n73_W_out, 
            c2_n74_W_out=> c2_n74_W_out, 
            c2_n75_W_out=> c2_n75_W_out, 
            c2_n76_W_out=> c2_n76_W_out, 
            c2_n77_W_out=> c2_n77_W_out, 
            c2_n78_W_out=> c2_n78_W_out, 
            c2_n79_W_out=> c2_n79_W_out, 
            c2_n80_W_out=> c2_n80_W_out, 
            c2_n81_W_out=> c2_n81_W_out, 
            c2_n82_W_out=> c2_n82_W_out, 
            c2_n83_W_out=> c2_n83_W_out, 
            c2_n84_W_out=> c2_n84_W_out, 
            c2_n85_W_out=> c2_n85_W_out, 
            c2_n86_W_out=> c2_n86_W_out, 
            c2_n87_W_out=> c2_n87_W_out, 
            c2_n88_W_out=> c2_n88_W_out, 
            c2_n89_W_out=> c2_n89_W_out, 
            c2_n90_W_out=> c2_n90_W_out, 
            c2_n91_W_out=> c2_n91_W_out, 
            c2_n92_W_out=> c2_n92_W_out, 
            c2_n93_W_out=> c2_n93_W_out, 
            c2_n94_W_out=> c2_n94_W_out, 
            c2_n95_W_out=> c2_n95_W_out, 
            c2_n96_W_out=> c2_n96_W_out, 
            c2_n97_W_out=> c2_n97_W_out, 
            c2_n98_W_out=> c2_n98_W_out, 
            c2_n99_W_out=> c2_n99_W_out
   );
            
camada3_inst_3: ENTITY work.camada3_ReLU_300neuron_8bits_100n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c3_IO_in, 
            c3_n0_W_in=> c2_n0_W_out,
            c3_n1_W_in=> c2_n1_W_out,
            c3_n2_W_in=> c2_n2_W_out,
            c3_n3_W_in=> c2_n3_W_out,
            c3_n4_W_in=> c2_n4_W_out,
            c3_n5_W_in=> c2_n5_W_out,
            c3_n6_W_in=> c2_n6_W_out,
            c3_n7_W_in=> c2_n7_W_out,
            c3_n8_W_in=> c2_n8_W_out,
            c3_n9_W_in=> c2_n9_W_out,
            c3_n10_W_in=> c2_n10_W_out,
            c3_n11_W_in=> c2_n11_W_out,
            c3_n12_W_in=> c2_n12_W_out,
            c3_n13_W_in=> c2_n13_W_out,
            c3_n14_W_in=> c2_n14_W_out,
            c3_n15_W_in=> c2_n15_W_out,
            c3_n16_W_in=> c2_n16_W_out,
            c3_n17_W_in=> c2_n17_W_out,
            c3_n18_W_in=> c2_n18_W_out,
            c3_n19_W_in=> c2_n19_W_out,
            c3_n20_W_in=> c2_n20_W_out,
            c3_n21_W_in=> c2_n21_W_out,
            c3_n22_W_in=> c2_n22_W_out,
            c3_n23_W_in=> c2_n23_W_out,
            c3_n24_W_in=> c2_n24_W_out,
            c3_n25_W_in=> c2_n25_W_out,
            c3_n26_W_in=> c2_n26_W_out,
            c3_n27_W_in=> c2_n27_W_out,
            c3_n28_W_in=> c2_n28_W_out,
            c3_n29_W_in=> c2_n29_W_out,
            c3_n30_W_in=> c2_n30_W_out,
            c3_n31_W_in=> c2_n31_W_out,
            c3_n32_W_in=> c2_n32_W_out,
            c3_n33_W_in=> c2_n33_W_out,
            c3_n34_W_in=> c2_n34_W_out,
            c3_n35_W_in=> c2_n35_W_out,
            c3_n36_W_in=> c2_n36_W_out,
            c3_n37_W_in=> c2_n37_W_out,
            c3_n38_W_in=> c2_n38_W_out,
            c3_n39_W_in=> c2_n39_W_out,
            c3_n40_W_in=> c2_n40_W_out,
            c3_n41_W_in=> c2_n41_W_out,
            c3_n42_W_in=> c2_n42_W_out,
            c3_n43_W_in=> c2_n43_W_out,
            c3_n44_W_in=> c2_n44_W_out,
            c3_n45_W_in=> c2_n45_W_out,
            c3_n46_W_in=> c2_n46_W_out,
            c3_n47_W_in=> c2_n47_W_out,
            c3_n48_W_in=> c2_n48_W_out,
            c3_n49_W_in=> c2_n49_W_out,
            c3_n50_W_in=> c2_n50_W_out,
            c3_n51_W_in=> c2_n51_W_out,
            c3_n52_W_in=> c2_n52_W_out,
            c3_n53_W_in=> c2_n53_W_out,
            c3_n54_W_in=> c2_n54_W_out,
            c3_n55_W_in=> c2_n55_W_out,
            c3_n56_W_in=> c2_n56_W_out,
            c3_n57_W_in=> c2_n57_W_out,
            c3_n58_W_in=> c2_n58_W_out,
            c3_n59_W_in=> c2_n59_W_out,
            c3_n60_W_in=> c2_n60_W_out,
            c3_n61_W_in=> c2_n61_W_out,
            c3_n62_W_in=> c2_n62_W_out,
            c3_n63_W_in=> c2_n63_W_out,
            c3_n64_W_in=> c2_n64_W_out,
            c3_n65_W_in=> c2_n65_W_out,
            c3_n66_W_in=> c2_n66_W_out,
            c3_n67_W_in=> c2_n67_W_out,
            c3_n68_W_in=> c2_n68_W_out,
            c3_n69_W_in=> c2_n69_W_out,
            c3_n70_W_in=> c2_n70_W_out,
            c3_n71_W_in=> c2_n71_W_out,
            c3_n72_W_in=> c2_n72_W_out,
            c3_n73_W_in=> c2_n73_W_out,
            c3_n74_W_in=> c2_n74_W_out,
            c3_n75_W_in=> c2_n75_W_out,
            c3_n76_W_in=> c2_n76_W_out,
            c3_n77_W_in=> c2_n77_W_out,
            c3_n78_W_in=> c2_n78_W_out,
            c3_n79_W_in=> c2_n79_W_out,
            c3_n80_W_in=> c2_n80_W_out,
            c3_n81_W_in=> c2_n81_W_out,
            c3_n82_W_in=> c2_n82_W_out,
            c3_n83_W_in=> c2_n83_W_out,
            c3_n84_W_in=> c2_n84_W_out,
            c3_n85_W_in=> c2_n85_W_out,
            c3_n86_W_in=> c2_n86_W_out,
            c3_n87_W_in=> c2_n87_W_out,
            c3_n88_W_in=> c2_n88_W_out,
            c3_n89_W_in=> c2_n89_W_out,
            c3_n90_W_in=> c2_n90_W_out,
            c3_n91_W_in=> c2_n91_W_out,
            c3_n92_W_in=> c2_n92_W_out,
            c3_n93_W_in=> c2_n93_W_out,
            c3_n94_W_in=> c2_n94_W_out,
            c3_n95_W_in=> c2_n95_W_out,
            c3_n96_W_in=> c2_n96_W_out,
            c3_n97_W_in=> c2_n97_W_out,
            c3_n98_W_in=> c2_n98_W_out,
            c3_n99_W_in=> c2_n99_W_out,
            c3_n100_W_in=> c1_n100_W_out,
            c3_n101_W_in=> c1_n101_W_out,
            c3_n102_W_in=> c1_n102_W_out,
            c3_n103_W_in=> c1_n103_W_out,
            c3_n104_W_in=> c1_n104_W_out,
            c3_n105_W_in=> c1_n105_W_out,
            c3_n106_W_in=> c1_n106_W_out,
            c3_n107_W_in=> c1_n107_W_out,
            c3_n108_W_in=> c1_n108_W_out,
            c3_n109_W_in=> c1_n109_W_out,
            c3_n110_W_in=> c1_n110_W_out,
            c3_n111_W_in=> c1_n111_W_out,
            c3_n112_W_in=> c1_n112_W_out,
            c3_n113_W_in=> c1_n113_W_out,
            c3_n114_W_in=> c1_n114_W_out,
            c3_n115_W_in=> c1_n115_W_out,
            c3_n116_W_in=> c1_n116_W_out,
            c3_n117_W_in=> c1_n117_W_out,
            c3_n118_W_in=> c1_n118_W_out,
            c3_n119_W_in=> c1_n119_W_out,
            c3_n120_W_in=> c1_n120_W_out,
            c3_n121_W_in=> c1_n121_W_out,
            c3_n122_W_in=> c1_n122_W_out,
            c3_n123_W_in=> c1_n123_W_out,
            c3_n124_W_in=> c1_n124_W_out,
            c3_n125_W_in=> c1_n125_W_out,
            c3_n126_W_in=> c1_n126_W_out,
            c3_n127_W_in=> c1_n127_W_out,
            c3_n128_W_in=> c1_n128_W_out,
            c3_n129_W_in=> c1_n129_W_out,
            c3_n130_W_in=> c1_n130_W_out,
            c3_n131_W_in=> c1_n131_W_out,
            c3_n132_W_in=> c1_n132_W_out,
            c3_n133_W_in=> c1_n133_W_out,
            c3_n134_W_in=> c1_n134_W_out,
            c3_n135_W_in=> c1_n135_W_out,
            c3_n136_W_in=> c1_n136_W_out,
            c3_n137_W_in=> c1_n137_W_out,
            c3_n138_W_in=> c1_n138_W_out,
            c3_n139_W_in=> c1_n139_W_out,
            c3_n140_W_in=> c1_n140_W_out,
            c3_n141_W_in=> c1_n141_W_out,
            c3_n142_W_in=> c1_n142_W_out,
            c3_n143_W_in=> c1_n143_W_out,
            c3_n144_W_in=> c1_n144_W_out,
            c3_n145_W_in=> c1_n145_W_out,
            c3_n146_W_in=> c1_n146_W_out,
            c3_n147_W_in=> c1_n147_W_out,
            c3_n148_W_in=> c1_n148_W_out,
            c3_n149_W_in=> c1_n149_W_out,
            c3_n150_W_in=> c1_n150_W_out,
            c3_n151_W_in=> c1_n151_W_out,
            c3_n152_W_in=> c1_n152_W_out,
            c3_n153_W_in=> c1_n153_W_out,
            c3_n154_W_in=> c1_n154_W_out,
            c3_n155_W_in=> c1_n155_W_out,
            c3_n156_W_in=> c1_n156_W_out,
            c3_n157_W_in=> c1_n157_W_out,
            c3_n158_W_in=> c1_n158_W_out,
            c3_n159_W_in=> c1_n159_W_out,
            c3_n160_W_in=> c1_n160_W_out,
            c3_n161_W_in=> c1_n161_W_out,
            c3_n162_W_in=> c1_n162_W_out,
            c3_n163_W_in=> c1_n163_W_out,
            c3_n164_W_in=> c1_n164_W_out,
            c3_n165_W_in=> c1_n165_W_out,
            c3_n166_W_in=> c1_n166_W_out,
            c3_n167_W_in=> c1_n167_W_out,
            c3_n168_W_in=> c1_n168_W_out,
            c3_n169_W_in=> c1_n169_W_out,
            c3_n170_W_in=> c1_n170_W_out,
            c3_n171_W_in=> c1_n171_W_out,
            c3_n172_W_in=> c1_n172_W_out,
            c3_n173_W_in=> c1_n173_W_out,
            c3_n174_W_in=> c1_n174_W_out,
            c3_n175_W_in=> c1_n175_W_out,
            c3_n176_W_in=> c1_n176_W_out,
            c3_n177_W_in=> c1_n177_W_out,
            c3_n178_W_in=> c1_n178_W_out,
            c3_n179_W_in=> c1_n179_W_out,
            c3_n180_W_in=> c1_n180_W_out,
            c3_n181_W_in=> c1_n181_W_out,
            c3_n182_W_in=> c1_n182_W_out,
            c3_n183_W_in=> c1_n183_W_out,
            c3_n184_W_in=> c1_n184_W_out,
            c3_n185_W_in=> c1_n185_W_out,
            c3_n186_W_in=> c1_n186_W_out,
            c3_n187_W_in=> c1_n187_W_out,
            c3_n188_W_in=> c1_n188_W_out,
            c3_n189_W_in=> c1_n189_W_out,
            c3_n190_W_in=> c1_n190_W_out,
            c3_n191_W_in=> c1_n191_W_out,
            c3_n192_W_in=> c1_n192_W_out,
            c3_n193_W_in=> c1_n193_W_out,
            c3_n194_W_in=> c1_n194_W_out,
            c3_n195_W_in=> c1_n195_W_out,
            c3_n196_W_in=> c1_n196_W_out,
            c3_n197_W_in=> c1_n197_W_out,
            c3_n198_W_in=> c1_n198_W_out,
            c3_n199_W_in=> c1_n199_W_out,
            c3_n200_W_in=> c1_n200_W_out,
            c3_n201_W_in=> c1_n201_W_out,
            c3_n202_W_in=> c1_n202_W_out,
            c3_n203_W_in=> c1_n203_W_out,
            c3_n204_W_in=> c1_n204_W_out,
            c3_n205_W_in=> c1_n205_W_out,
            c3_n206_W_in=> c1_n206_W_out,
            c3_n207_W_in=> c1_n207_W_out,
            c3_n208_W_in=> c1_n208_W_out,
            c3_n209_W_in=> c1_n209_W_out,
            c3_n210_W_in=> c1_n210_W_out,
            c3_n211_W_in=> c1_n211_W_out,
            c3_n212_W_in=> c1_n212_W_out,
            c3_n213_W_in=> c1_n213_W_out,
            c3_n214_W_in=> c1_n214_W_out,
            c3_n215_W_in=> c1_n215_W_out,
            c3_n216_W_in=> c1_n216_W_out,
            c3_n217_W_in=> c1_n217_W_out,
            c3_n218_W_in=> c1_n218_W_out,
            c3_n219_W_in=> c1_n219_W_out,
            c3_n220_W_in=> c1_n220_W_out,
            c3_n221_W_in=> c1_n221_W_out,
            c3_n222_W_in=> c1_n222_W_out,
            c3_n223_W_in=> c1_n223_W_out,
            c3_n224_W_in=> c1_n224_W_out,
            c3_n225_W_in=> c1_n225_W_out,
            c3_n226_W_in=> c1_n226_W_out,
            c3_n227_W_in=> c1_n227_W_out,
            c3_n228_W_in=> c1_n228_W_out,
            c3_n229_W_in=> c1_n229_W_out,
            c3_n230_W_in=> c1_n230_W_out,
            c3_n231_W_in=> c1_n231_W_out,
            c3_n232_W_in=> c1_n232_W_out,
            c3_n233_W_in=> c1_n233_W_out,
            c3_n234_W_in=> c1_n234_W_out,
            c3_n235_W_in=> c1_n235_W_out,
            c3_n236_W_in=> c1_n236_W_out,
            c3_n237_W_in=> c1_n237_W_out,
            c3_n238_W_in=> c1_n238_W_out,
            c3_n239_W_in=> c1_n239_W_out,
            c3_n240_W_in=> c1_n240_W_out,
            c3_n241_W_in=> c1_n241_W_out,
            c3_n242_W_in=> c1_n242_W_out,
            c3_n243_W_in=> c1_n243_W_out,
            c3_n244_W_in=> c1_n244_W_out,
            c3_n245_W_in=> c1_n245_W_out,
            c3_n246_W_in=> c1_n246_W_out,
            c3_n247_W_in=> c1_n247_W_out,
            c3_n248_W_in=> c1_n248_W_out,
            c3_n249_W_in=> c1_n249_W_out,
            c3_n250_W_in=> c1_n250_W_out,
            c3_n251_W_in=> c1_n251_W_out,
            c3_n252_W_in=> c1_n252_W_out,
            c3_n253_W_in=> c1_n253_W_out,
            c3_n254_W_in=> c1_n254_W_out,
            c3_n255_W_in=> c1_n255_W_out,
            c3_n256_W_in=> c1_n256_W_out,
            c3_n257_W_in=> c1_n257_W_out,
            c3_n258_W_in=> c1_n258_W_out,
            c3_n259_W_in=> c1_n259_W_out,
            c3_n260_W_in=> c1_n260_W_out,
            c3_n261_W_in=> c1_n261_W_out,
            c3_n262_W_in=> c1_n262_W_out,
            c3_n263_W_in=> c1_n263_W_out,
            c3_n264_W_in=> c1_n264_W_out,
            c3_n265_W_in=> c1_n265_W_out,
            c3_n266_W_in=> c1_n266_W_out,
            c3_n267_W_in=> c1_n267_W_out,
            c3_n268_W_in=> c1_n268_W_out,
            c3_n269_W_in=> c1_n269_W_out,
            c3_n270_W_in=> c1_n270_W_out,
            c3_n271_W_in=> c1_n271_W_out,
            c3_n272_W_in=> c1_n272_W_out,
            c3_n273_W_in=> c1_n273_W_out,
            c3_n274_W_in=> c1_n274_W_out,
            c3_n275_W_in=> c1_n275_W_out,
            c3_n276_W_in=> c1_n276_W_out,
            c3_n277_W_in=> c1_n277_W_out,
            c3_n278_W_in=> c1_n278_W_out,
            c3_n279_W_in=> c1_n279_W_out,
            c3_n280_W_in=> c1_n280_W_out,
            c3_n281_W_in=> c1_n281_W_out,
            c3_n282_W_in=> c1_n282_W_out,
            c3_n283_W_in=> c1_n283_W_out,
            c3_n284_W_in=> c1_n284_W_out,
            c3_n285_W_in=> c1_n285_W_out,
            c3_n286_W_in=> c1_n286_W_out,
            c3_n287_W_in=> c1_n287_W_out,
            c3_n288_W_in=> c1_n288_W_out,
            c3_n289_W_in=> c1_n289_W_out,
            c3_n290_W_in=> c1_n290_W_out,
            c3_n291_W_in=> c1_n291_W_out,
            c3_n292_W_in=> c1_n292_W_out,
            c3_n293_W_in=> c1_n293_W_out,
            c3_n294_W_in=> c1_n294_W_out,
            c3_n295_W_in=> c1_n295_W_out,
            c3_n296_W_in=> c1_n296_W_out,
            c3_n297_W_in=> c1_n297_W_out,
            c3_n298_W_in=> c1_n298_W_out,
            c3_n299_W_in=> c1_n299_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c3_n0_IO_out=> c3_n0_IO_out, 
            c3_n1_IO_out=> c3_n1_IO_out, 
            c3_n2_IO_out=> c3_n2_IO_out, 
            c3_n3_IO_out=> c3_n3_IO_out, 
            c3_n4_IO_out=> c3_n4_IO_out, 
            c3_n5_IO_out=> c3_n5_IO_out, 
            c3_n6_IO_out=> c3_n6_IO_out, 
            c3_n7_IO_out=> c3_n7_IO_out, 
            c3_n8_IO_out=> c3_n8_IO_out, 
            c3_n9_IO_out=> c3_n9_IO_out, 
            c3_n10_IO_out=> c3_n10_IO_out, 
            c3_n11_IO_out=> c3_n11_IO_out, 
            c3_n12_IO_out=> c3_n12_IO_out, 
            c3_n13_IO_out=> c3_n13_IO_out, 
            c3_n14_IO_out=> c3_n14_IO_out, 
            c3_n15_IO_out=> c3_n15_IO_out, 
            c3_n16_IO_out=> c3_n16_IO_out, 
            c3_n17_IO_out=> c3_n17_IO_out, 
            c3_n18_IO_out=> c3_n18_IO_out, 
            c3_n19_IO_out=> c3_n19_IO_out, 
            c3_n20_IO_out=> c3_n20_IO_out, 
            c3_n21_IO_out=> c3_n21_IO_out, 
            c3_n22_IO_out=> c3_n22_IO_out, 
            c3_n23_IO_out=> c3_n23_IO_out, 
            c3_n24_IO_out=> c3_n24_IO_out, 
            c3_n25_IO_out=> c3_n25_IO_out, 
            c3_n26_IO_out=> c3_n26_IO_out, 
            c3_n27_IO_out=> c3_n27_IO_out, 
            c3_n28_IO_out=> c3_n28_IO_out, 
            c3_n29_IO_out=> c3_n29_IO_out, 
            c3_n30_IO_out=> c3_n30_IO_out, 
            c3_n31_IO_out=> c3_n31_IO_out, 
            c3_n32_IO_out=> c3_n32_IO_out, 
            c3_n33_IO_out=> c3_n33_IO_out, 
            c3_n34_IO_out=> c3_n34_IO_out, 
            c3_n35_IO_out=> c3_n35_IO_out, 
            c3_n36_IO_out=> c3_n36_IO_out, 
            c3_n37_IO_out=> c3_n37_IO_out, 
            c3_n38_IO_out=> c3_n38_IO_out, 
            c3_n39_IO_out=> c3_n39_IO_out, 
            c3_n40_IO_out=> c3_n40_IO_out, 
            c3_n41_IO_out=> c3_n41_IO_out, 
            c3_n42_IO_out=> c3_n42_IO_out, 
            c3_n43_IO_out=> c3_n43_IO_out, 
            c3_n44_IO_out=> c3_n44_IO_out, 
            c3_n45_IO_out=> c3_n45_IO_out, 
            c3_n46_IO_out=> c3_n46_IO_out, 
            c3_n47_IO_out=> c3_n47_IO_out, 
            c3_n48_IO_out=> c3_n48_IO_out, 
            c3_n49_IO_out=> c3_n49_IO_out, 
            c3_n50_IO_out=> c3_n50_IO_out, 
            c3_n51_IO_out=> c3_n51_IO_out, 
            c3_n52_IO_out=> c3_n52_IO_out, 
            c3_n53_IO_out=> c3_n53_IO_out, 
            c3_n54_IO_out=> c3_n54_IO_out, 
            c3_n55_IO_out=> c3_n55_IO_out, 
            c3_n56_IO_out=> c3_n56_IO_out, 
            c3_n57_IO_out=> c3_n57_IO_out, 
            c3_n58_IO_out=> c3_n58_IO_out, 
            c3_n59_IO_out=> c3_n59_IO_out, 
            c3_n60_IO_out=> c3_n60_IO_out, 
            c3_n61_IO_out=> c3_n61_IO_out, 
            c3_n62_IO_out=> c3_n62_IO_out, 
            c3_n63_IO_out=> c3_n63_IO_out, 
            c3_n64_IO_out=> c3_n64_IO_out, 
            c3_n65_IO_out=> c3_n65_IO_out, 
            c3_n66_IO_out=> c3_n66_IO_out, 
            c3_n67_IO_out=> c3_n67_IO_out, 
            c3_n68_IO_out=> c3_n68_IO_out, 
            c3_n69_IO_out=> c3_n69_IO_out, 
            c3_n70_IO_out=> c3_n70_IO_out, 
            c3_n71_IO_out=> c3_n71_IO_out, 
            c3_n72_IO_out=> c3_n72_IO_out, 
            c3_n73_IO_out=> c3_n73_IO_out, 
            c3_n74_IO_out=> c3_n74_IO_out, 
            c3_n75_IO_out=> c3_n75_IO_out, 
            c3_n76_IO_out=> c3_n76_IO_out, 
            c3_n77_IO_out=> c3_n77_IO_out, 
            c3_n78_IO_out=> c3_n78_IO_out, 
            c3_n79_IO_out=> c3_n79_IO_out, 
            c3_n80_IO_out=> c3_n80_IO_out, 
            c3_n81_IO_out=> c3_n81_IO_out, 
            c3_n82_IO_out=> c3_n82_IO_out, 
            c3_n83_IO_out=> c3_n83_IO_out, 
            c3_n84_IO_out=> c3_n84_IO_out, 
            c3_n85_IO_out=> c3_n85_IO_out, 
            c3_n86_IO_out=> c3_n86_IO_out, 
            c3_n87_IO_out=> c3_n87_IO_out, 
            c3_n88_IO_out=> c3_n88_IO_out, 
            c3_n89_IO_out=> c3_n89_IO_out, 
            c3_n90_IO_out=> c3_n90_IO_out, 
            c3_n91_IO_out=> c3_n91_IO_out, 
            c3_n92_IO_out=> c3_n92_IO_out, 
            c3_n93_IO_out=> c3_n93_IO_out, 
            c3_n94_IO_out=> c3_n94_IO_out, 
            c3_n95_IO_out=> c3_n95_IO_out, 
            c3_n96_IO_out=> c3_n96_IO_out, 
            c3_n97_IO_out=> c3_n97_IO_out, 
            c3_n98_IO_out=> c3_n98_IO_out, 
            c3_n99_IO_out=> c3_n99_IO_out, 
            c3_n100_IO_out=> c3_n100_IO_out, 
            c3_n101_IO_out=> c3_n101_IO_out, 
            c3_n102_IO_out=> c3_n102_IO_out, 
            c3_n103_IO_out=> c3_n103_IO_out, 
            c3_n104_IO_out=> c3_n104_IO_out, 
            c3_n105_IO_out=> c3_n105_IO_out, 
            c3_n106_IO_out=> c3_n106_IO_out, 
            c3_n107_IO_out=> c3_n107_IO_out, 
            c3_n108_IO_out=> c3_n108_IO_out, 
            c3_n109_IO_out=> c3_n109_IO_out, 
            c3_n110_IO_out=> c3_n110_IO_out, 
            c3_n111_IO_out=> c3_n111_IO_out, 
            c3_n112_IO_out=> c3_n112_IO_out, 
            c3_n113_IO_out=> c3_n113_IO_out, 
            c3_n114_IO_out=> c3_n114_IO_out, 
            c3_n115_IO_out=> c3_n115_IO_out, 
            c3_n116_IO_out=> c3_n116_IO_out, 
            c3_n117_IO_out=> c3_n117_IO_out, 
            c3_n118_IO_out=> c3_n118_IO_out, 
            c3_n119_IO_out=> c3_n119_IO_out, 
            c3_n120_IO_out=> c3_n120_IO_out, 
            c3_n121_IO_out=> c3_n121_IO_out, 
            c3_n122_IO_out=> c3_n122_IO_out, 
            c3_n123_IO_out=> c3_n123_IO_out, 
            c3_n124_IO_out=> c3_n124_IO_out, 
            c3_n125_IO_out=> c3_n125_IO_out, 
            c3_n126_IO_out=> c3_n126_IO_out, 
            c3_n127_IO_out=> c3_n127_IO_out, 
            c3_n128_IO_out=> c3_n128_IO_out, 
            c3_n129_IO_out=> c3_n129_IO_out, 
            c3_n130_IO_out=> c3_n130_IO_out, 
            c3_n131_IO_out=> c3_n131_IO_out, 
            c3_n132_IO_out=> c3_n132_IO_out, 
            c3_n133_IO_out=> c3_n133_IO_out, 
            c3_n134_IO_out=> c3_n134_IO_out, 
            c3_n135_IO_out=> c3_n135_IO_out, 
            c3_n136_IO_out=> c3_n136_IO_out, 
            c3_n137_IO_out=> c3_n137_IO_out, 
            c3_n138_IO_out=> c3_n138_IO_out, 
            c3_n139_IO_out=> c3_n139_IO_out, 
            c3_n140_IO_out=> c3_n140_IO_out, 
            c3_n141_IO_out=> c3_n141_IO_out, 
            c3_n142_IO_out=> c3_n142_IO_out, 
            c3_n143_IO_out=> c3_n143_IO_out, 
            c3_n144_IO_out=> c3_n144_IO_out, 
            c3_n145_IO_out=> c3_n145_IO_out, 
            c3_n146_IO_out=> c3_n146_IO_out, 
            c3_n147_IO_out=> c3_n147_IO_out, 
            c3_n148_IO_out=> c3_n148_IO_out, 
            c3_n149_IO_out=> c3_n149_IO_out, 
            c3_n150_IO_out=> c3_n150_IO_out, 
            c3_n151_IO_out=> c3_n151_IO_out, 
            c3_n152_IO_out=> c3_n152_IO_out, 
            c3_n153_IO_out=> c3_n153_IO_out, 
            c3_n154_IO_out=> c3_n154_IO_out, 
            c3_n155_IO_out=> c3_n155_IO_out, 
            c3_n156_IO_out=> c3_n156_IO_out, 
            c3_n157_IO_out=> c3_n157_IO_out, 
            c3_n158_IO_out=> c3_n158_IO_out, 
            c3_n159_IO_out=> c3_n159_IO_out, 
            c3_n160_IO_out=> c3_n160_IO_out, 
            c3_n161_IO_out=> c3_n161_IO_out, 
            c3_n162_IO_out=> c3_n162_IO_out, 
            c3_n163_IO_out=> c3_n163_IO_out, 
            c3_n164_IO_out=> c3_n164_IO_out, 
            c3_n165_IO_out=> c3_n165_IO_out, 
            c3_n166_IO_out=> c3_n166_IO_out, 
            c3_n167_IO_out=> c3_n167_IO_out, 
            c3_n168_IO_out=> c3_n168_IO_out, 
            c3_n169_IO_out=> c3_n169_IO_out, 
            c3_n170_IO_out=> c3_n170_IO_out, 
            c3_n171_IO_out=> c3_n171_IO_out, 
            c3_n172_IO_out=> c3_n172_IO_out, 
            c3_n173_IO_out=> c3_n173_IO_out, 
            c3_n174_IO_out=> c3_n174_IO_out, 
            c3_n175_IO_out=> c3_n175_IO_out, 
            c3_n176_IO_out=> c3_n176_IO_out, 
            c3_n177_IO_out=> c3_n177_IO_out, 
            c3_n178_IO_out=> c3_n178_IO_out, 
            c3_n179_IO_out=> c3_n179_IO_out, 
            c3_n180_IO_out=> c3_n180_IO_out, 
            c3_n181_IO_out=> c3_n181_IO_out, 
            c3_n182_IO_out=> c3_n182_IO_out, 
            c3_n183_IO_out=> c3_n183_IO_out, 
            c3_n184_IO_out=> c3_n184_IO_out, 
            c3_n185_IO_out=> c3_n185_IO_out, 
            c3_n186_IO_out=> c3_n186_IO_out, 
            c3_n187_IO_out=> c3_n187_IO_out, 
            c3_n188_IO_out=> c3_n188_IO_out, 
            c3_n189_IO_out=> c3_n189_IO_out, 
            c3_n190_IO_out=> c3_n190_IO_out, 
            c3_n191_IO_out=> c3_n191_IO_out, 
            c3_n192_IO_out=> c3_n192_IO_out, 
            c3_n193_IO_out=> c3_n193_IO_out, 
            c3_n194_IO_out=> c3_n194_IO_out, 
            c3_n195_IO_out=> c3_n195_IO_out, 
            c3_n196_IO_out=> c3_n196_IO_out, 
            c3_n197_IO_out=> c3_n197_IO_out, 
            c3_n198_IO_out=> c3_n198_IO_out, 
            c3_n199_IO_out=> c3_n199_IO_out, 
            c3_n200_IO_out=> c3_n200_IO_out, 
            c3_n201_IO_out=> c3_n201_IO_out, 
            c3_n202_IO_out=> c3_n202_IO_out, 
            c3_n203_IO_out=> c3_n203_IO_out, 
            c3_n204_IO_out=> c3_n204_IO_out, 
            c3_n205_IO_out=> c3_n205_IO_out, 
            c3_n206_IO_out=> c3_n206_IO_out, 
            c3_n207_IO_out=> c3_n207_IO_out, 
            c3_n208_IO_out=> c3_n208_IO_out, 
            c3_n209_IO_out=> c3_n209_IO_out, 
            c3_n210_IO_out=> c3_n210_IO_out, 
            c3_n211_IO_out=> c3_n211_IO_out, 
            c3_n212_IO_out=> c3_n212_IO_out, 
            c3_n213_IO_out=> c3_n213_IO_out, 
            c3_n214_IO_out=> c3_n214_IO_out, 
            c3_n215_IO_out=> c3_n215_IO_out, 
            c3_n216_IO_out=> c3_n216_IO_out, 
            c3_n217_IO_out=> c3_n217_IO_out, 
            c3_n218_IO_out=> c3_n218_IO_out, 
            c3_n219_IO_out=> c3_n219_IO_out, 
            c3_n220_IO_out=> c3_n220_IO_out, 
            c3_n221_IO_out=> c3_n221_IO_out, 
            c3_n222_IO_out=> c3_n222_IO_out, 
            c3_n223_IO_out=> c3_n223_IO_out, 
            c3_n224_IO_out=> c3_n224_IO_out, 
            c3_n225_IO_out=> c3_n225_IO_out, 
            c3_n226_IO_out=> c3_n226_IO_out, 
            c3_n227_IO_out=> c3_n227_IO_out, 
            c3_n228_IO_out=> c3_n228_IO_out, 
            c3_n229_IO_out=> c3_n229_IO_out, 
            c3_n230_IO_out=> c3_n230_IO_out, 
            c3_n231_IO_out=> c3_n231_IO_out, 
            c3_n232_IO_out=> c3_n232_IO_out, 
            c3_n233_IO_out=> c3_n233_IO_out, 
            c3_n234_IO_out=> c3_n234_IO_out, 
            c3_n235_IO_out=> c3_n235_IO_out, 
            c3_n236_IO_out=> c3_n236_IO_out, 
            c3_n237_IO_out=> c3_n237_IO_out, 
            c3_n238_IO_out=> c3_n238_IO_out, 
            c3_n239_IO_out=> c3_n239_IO_out, 
            c3_n240_IO_out=> c3_n240_IO_out, 
            c3_n241_IO_out=> c3_n241_IO_out, 
            c3_n242_IO_out=> c3_n242_IO_out, 
            c3_n243_IO_out=> c3_n243_IO_out, 
            c3_n244_IO_out=> c3_n244_IO_out, 
            c3_n245_IO_out=> c3_n245_IO_out, 
            c3_n246_IO_out=> c3_n246_IO_out, 
            c3_n247_IO_out=> c3_n247_IO_out, 
            c3_n248_IO_out=> c3_n248_IO_out, 
            c3_n249_IO_out=> c3_n249_IO_out, 
            c3_n250_IO_out=> c3_n250_IO_out, 
            c3_n251_IO_out=> c3_n251_IO_out, 
            c3_n252_IO_out=> c3_n252_IO_out, 
            c3_n253_IO_out=> c3_n253_IO_out, 
            c3_n254_IO_out=> c3_n254_IO_out, 
            c3_n255_IO_out=> c3_n255_IO_out, 
            c3_n256_IO_out=> c3_n256_IO_out, 
            c3_n257_IO_out=> c3_n257_IO_out, 
            c3_n258_IO_out=> c3_n258_IO_out, 
            c3_n259_IO_out=> c3_n259_IO_out, 
            c3_n260_IO_out=> c3_n260_IO_out, 
            c3_n261_IO_out=> c3_n261_IO_out, 
            c3_n262_IO_out=> c3_n262_IO_out, 
            c3_n263_IO_out=> c3_n263_IO_out, 
            c3_n264_IO_out=> c3_n264_IO_out, 
            c3_n265_IO_out=> c3_n265_IO_out, 
            c3_n266_IO_out=> c3_n266_IO_out, 
            c3_n267_IO_out=> c3_n267_IO_out, 
            c3_n268_IO_out=> c3_n268_IO_out, 
            c3_n269_IO_out=> c3_n269_IO_out, 
            c3_n270_IO_out=> c3_n270_IO_out, 
            c3_n271_IO_out=> c3_n271_IO_out, 
            c3_n272_IO_out=> c3_n272_IO_out, 
            c3_n273_IO_out=> c3_n273_IO_out, 
            c3_n274_IO_out=> c3_n274_IO_out, 
            c3_n275_IO_out=> c3_n275_IO_out, 
            c3_n276_IO_out=> c3_n276_IO_out, 
            c3_n277_IO_out=> c3_n277_IO_out, 
            c3_n278_IO_out=> c3_n278_IO_out, 
            c3_n279_IO_out=> c3_n279_IO_out, 
            c3_n280_IO_out=> c3_n280_IO_out, 
            c3_n281_IO_out=> c3_n281_IO_out, 
            c3_n282_IO_out=> c3_n282_IO_out, 
            c3_n283_IO_out=> c3_n283_IO_out, 
            c3_n284_IO_out=> c3_n284_IO_out, 
            c3_n285_IO_out=> c3_n285_IO_out, 
            c3_n286_IO_out=> c3_n286_IO_out, 
            c3_n287_IO_out=> c3_n287_IO_out, 
            c3_n288_IO_out=> c3_n288_IO_out, 
            c3_n289_IO_out=> c3_n289_IO_out, 
            c3_n290_IO_out=> c3_n290_IO_out, 
            c3_n291_IO_out=> c3_n291_IO_out, 
            c3_n292_IO_out=> c3_n292_IO_out, 
            c3_n293_IO_out=> c3_n293_IO_out, 
            c3_n294_IO_out=> c3_n294_IO_out, 
            c3_n295_IO_out=> c3_n295_IO_out, 
            c3_n296_IO_out=> c3_n296_IO_out, 
            c3_n297_IO_out=> c3_n297_IO_out, 
            c3_n298_IO_out=> c3_n298_IO_out, 
            c3_n299_IO_out=> c3_n299_IO_out, 
            -- ['OUT']['manual'] 
            c3_n0_W_out=> c3_n0_W_out, 
            c3_n1_W_out=> c3_n1_W_out, 
            c3_n2_W_out=> c3_n2_W_out, 
            c3_n3_W_out=> c3_n3_W_out, 
            c3_n4_W_out=> c3_n4_W_out, 
            c3_n5_W_out=> c3_n5_W_out, 
            c3_n6_W_out=> c3_n6_W_out, 
            c3_n7_W_out=> c3_n7_W_out, 
            c3_n8_W_out=> c3_n8_W_out, 
            c3_n9_W_out=> c3_n9_W_out, 
            c3_n10_W_out=> c3_n10_W_out, 
            c3_n11_W_out=> c3_n11_W_out, 
            c3_n12_W_out=> c3_n12_W_out, 
            c3_n13_W_out=> c3_n13_W_out, 
            c3_n14_W_out=> c3_n14_W_out, 
            c3_n15_W_out=> c3_n15_W_out, 
            c3_n16_W_out=> c3_n16_W_out, 
            c3_n17_W_out=> c3_n17_W_out, 
            c3_n18_W_out=> c3_n18_W_out, 
            c3_n19_W_out=> c3_n19_W_out, 
            c3_n20_W_out=> c3_n20_W_out, 
            c3_n21_W_out=> c3_n21_W_out, 
            c3_n22_W_out=> c3_n22_W_out, 
            c3_n23_W_out=> c3_n23_W_out, 
            c3_n24_W_out=> c3_n24_W_out, 
            c3_n25_W_out=> c3_n25_W_out, 
            c3_n26_W_out=> c3_n26_W_out, 
            c3_n27_W_out=> c3_n27_W_out, 
            c3_n28_W_out=> c3_n28_W_out, 
            c3_n29_W_out=> c3_n29_W_out, 
            c3_n30_W_out=> c3_n30_W_out, 
            c3_n31_W_out=> c3_n31_W_out, 
            c3_n32_W_out=> c3_n32_W_out, 
            c3_n33_W_out=> c3_n33_W_out, 
            c3_n34_W_out=> c3_n34_W_out, 
            c3_n35_W_out=> c3_n35_W_out, 
            c3_n36_W_out=> c3_n36_W_out, 
            c3_n37_W_out=> c3_n37_W_out, 
            c3_n38_W_out=> c3_n38_W_out, 
            c3_n39_W_out=> c3_n39_W_out, 
            c3_n40_W_out=> c3_n40_W_out, 
            c3_n41_W_out=> c3_n41_W_out, 
            c3_n42_W_out=> c3_n42_W_out, 
            c3_n43_W_out=> c3_n43_W_out, 
            c3_n44_W_out=> c3_n44_W_out, 
            c3_n45_W_out=> c3_n45_W_out, 
            c3_n46_W_out=> c3_n46_W_out, 
            c3_n47_W_out=> c3_n47_W_out, 
            c3_n48_W_out=> c3_n48_W_out, 
            c3_n49_W_out=> c3_n49_W_out, 
            c3_n50_W_out=> c3_n50_W_out, 
            c3_n51_W_out=> c3_n51_W_out, 
            c3_n52_W_out=> c3_n52_W_out, 
            c3_n53_W_out=> c3_n53_W_out, 
            c3_n54_W_out=> c3_n54_W_out, 
            c3_n55_W_out=> c3_n55_W_out, 
            c3_n56_W_out=> c3_n56_W_out, 
            c3_n57_W_out=> c3_n57_W_out, 
            c3_n58_W_out=> c3_n58_W_out, 
            c3_n59_W_out=> c3_n59_W_out, 
            c3_n60_W_out=> c3_n60_W_out, 
            c3_n61_W_out=> c3_n61_W_out, 
            c3_n62_W_out=> c3_n62_W_out, 
            c3_n63_W_out=> c3_n63_W_out, 
            c3_n64_W_out=> c3_n64_W_out, 
            c3_n65_W_out=> c3_n65_W_out, 
            c3_n66_W_out=> c3_n66_W_out, 
            c3_n67_W_out=> c3_n67_W_out, 
            c3_n68_W_out=> c3_n68_W_out, 
            c3_n69_W_out=> c3_n69_W_out, 
            c3_n70_W_out=> c3_n70_W_out, 
            c3_n71_W_out=> c3_n71_W_out, 
            c3_n72_W_out=> c3_n72_W_out, 
            c3_n73_W_out=> c3_n73_W_out, 
            c3_n74_W_out=> c3_n74_W_out, 
            c3_n75_W_out=> c3_n75_W_out, 
            c3_n76_W_out=> c3_n76_W_out, 
            c3_n77_W_out=> c3_n77_W_out, 
            c3_n78_W_out=> c3_n78_W_out, 
            c3_n79_W_out=> c3_n79_W_out, 
            c3_n80_W_out=> c3_n80_W_out, 
            c3_n81_W_out=> c3_n81_W_out, 
            c3_n82_W_out=> c3_n82_W_out, 
            c3_n83_W_out=> c3_n83_W_out, 
            c3_n84_W_out=> c3_n84_W_out, 
            c3_n85_W_out=> c3_n85_W_out, 
            c3_n86_W_out=> c3_n86_W_out, 
            c3_n87_W_out=> c3_n87_W_out, 
            c3_n88_W_out=> c3_n88_W_out, 
            c3_n89_W_out=> c3_n89_W_out, 
            c3_n90_W_out=> c3_n90_W_out, 
            c3_n91_W_out=> c3_n91_W_out, 
            c3_n92_W_out=> c3_n92_W_out, 
            c3_n93_W_out=> c3_n93_W_out, 
            c3_n94_W_out=> c3_n94_W_out, 
            c3_n95_W_out=> c3_n95_W_out, 
            c3_n96_W_out=> c3_n96_W_out, 
            c3_n97_W_out=> c3_n97_W_out, 
            c3_n98_W_out=> c3_n98_W_out, 
            c3_n99_W_out=> c3_n99_W_out, 
            c3_n100_W_out=> c3_n100_W_out, 
            c3_n101_W_out=> c3_n101_W_out, 
            c3_n102_W_out=> c3_n102_W_out, 
            c3_n103_W_out=> c3_n103_W_out, 
            c3_n104_W_out=> c3_n104_W_out, 
            c3_n105_W_out=> c3_n105_W_out, 
            c3_n106_W_out=> c3_n106_W_out, 
            c3_n107_W_out=> c3_n107_W_out, 
            c3_n108_W_out=> c3_n108_W_out, 
            c3_n109_W_out=> c3_n109_W_out, 
            c3_n110_W_out=> c3_n110_W_out, 
            c3_n111_W_out=> c3_n111_W_out, 
            c3_n112_W_out=> c3_n112_W_out, 
            c3_n113_W_out=> c3_n113_W_out, 
            c3_n114_W_out=> c3_n114_W_out, 
            c3_n115_W_out=> c3_n115_W_out, 
            c3_n116_W_out=> c3_n116_W_out, 
            c3_n117_W_out=> c3_n117_W_out, 
            c3_n118_W_out=> c3_n118_W_out, 
            c3_n119_W_out=> c3_n119_W_out, 
            c3_n120_W_out=> c3_n120_W_out, 
            c3_n121_W_out=> c3_n121_W_out, 
            c3_n122_W_out=> c3_n122_W_out, 
            c3_n123_W_out=> c3_n123_W_out, 
            c3_n124_W_out=> c3_n124_W_out, 
            c3_n125_W_out=> c3_n125_W_out, 
            c3_n126_W_out=> c3_n126_W_out, 
            c3_n127_W_out=> c3_n127_W_out, 
            c3_n128_W_out=> c3_n128_W_out, 
            c3_n129_W_out=> c3_n129_W_out, 
            c3_n130_W_out=> c3_n130_W_out, 
            c3_n131_W_out=> c3_n131_W_out, 
            c3_n132_W_out=> c3_n132_W_out, 
            c3_n133_W_out=> c3_n133_W_out, 
            c3_n134_W_out=> c3_n134_W_out, 
            c3_n135_W_out=> c3_n135_W_out, 
            c3_n136_W_out=> c3_n136_W_out, 
            c3_n137_W_out=> c3_n137_W_out, 
            c3_n138_W_out=> c3_n138_W_out, 
            c3_n139_W_out=> c3_n139_W_out, 
            c3_n140_W_out=> c3_n140_W_out, 
            c3_n141_W_out=> c3_n141_W_out, 
            c3_n142_W_out=> c3_n142_W_out, 
            c3_n143_W_out=> c3_n143_W_out, 
            c3_n144_W_out=> c3_n144_W_out, 
            c3_n145_W_out=> c3_n145_W_out, 
            c3_n146_W_out=> c3_n146_W_out, 
            c3_n147_W_out=> c3_n147_W_out, 
            c3_n148_W_out=> c3_n148_W_out, 
            c3_n149_W_out=> c3_n149_W_out, 
            c3_n150_W_out=> c3_n150_W_out, 
            c3_n151_W_out=> c3_n151_W_out, 
            c3_n152_W_out=> c3_n152_W_out, 
            c3_n153_W_out=> c3_n153_W_out, 
            c3_n154_W_out=> c3_n154_W_out, 
            c3_n155_W_out=> c3_n155_W_out, 
            c3_n156_W_out=> c3_n156_W_out, 
            c3_n157_W_out=> c3_n157_W_out, 
            c3_n158_W_out=> c3_n158_W_out, 
            c3_n159_W_out=> c3_n159_W_out, 
            c3_n160_W_out=> c3_n160_W_out, 
            c3_n161_W_out=> c3_n161_W_out, 
            c3_n162_W_out=> c3_n162_W_out, 
            c3_n163_W_out=> c3_n163_W_out, 
            c3_n164_W_out=> c3_n164_W_out, 
            c3_n165_W_out=> c3_n165_W_out, 
            c3_n166_W_out=> c3_n166_W_out, 
            c3_n167_W_out=> c3_n167_W_out, 
            c3_n168_W_out=> c3_n168_W_out, 
            c3_n169_W_out=> c3_n169_W_out, 
            c3_n170_W_out=> c3_n170_W_out, 
            c3_n171_W_out=> c3_n171_W_out, 
            c3_n172_W_out=> c3_n172_W_out, 
            c3_n173_W_out=> c3_n173_W_out, 
            c3_n174_W_out=> c3_n174_W_out, 
            c3_n175_W_out=> c3_n175_W_out, 
            c3_n176_W_out=> c3_n176_W_out, 
            c3_n177_W_out=> c3_n177_W_out, 
            c3_n178_W_out=> c3_n178_W_out, 
            c3_n179_W_out=> c3_n179_W_out, 
            c3_n180_W_out=> c3_n180_W_out, 
            c3_n181_W_out=> c3_n181_W_out, 
            c3_n182_W_out=> c3_n182_W_out, 
            c3_n183_W_out=> c3_n183_W_out, 
            c3_n184_W_out=> c3_n184_W_out, 
            c3_n185_W_out=> c3_n185_W_out, 
            c3_n186_W_out=> c3_n186_W_out, 
            c3_n187_W_out=> c3_n187_W_out, 
            c3_n188_W_out=> c3_n188_W_out, 
            c3_n189_W_out=> c3_n189_W_out, 
            c3_n190_W_out=> c3_n190_W_out, 
            c3_n191_W_out=> c3_n191_W_out, 
            c3_n192_W_out=> c3_n192_W_out, 
            c3_n193_W_out=> c3_n193_W_out, 
            c3_n194_W_out=> c3_n194_W_out, 
            c3_n195_W_out=> c3_n195_W_out, 
            c3_n196_W_out=> c3_n196_W_out, 
            c3_n197_W_out=> c3_n197_W_out, 
            c3_n198_W_out=> c3_n198_W_out, 
            c3_n199_W_out=> c3_n199_W_out, 
            c3_n200_W_out=> c3_n200_W_out, 
            c3_n201_W_out=> c3_n201_W_out, 
            c3_n202_W_out=> c3_n202_W_out, 
            c3_n203_W_out=> c3_n203_W_out, 
            c3_n204_W_out=> c3_n204_W_out, 
            c3_n205_W_out=> c3_n205_W_out, 
            c3_n206_W_out=> c3_n206_W_out, 
            c3_n207_W_out=> c3_n207_W_out, 
            c3_n208_W_out=> c3_n208_W_out, 
            c3_n209_W_out=> c3_n209_W_out, 
            c3_n210_W_out=> c3_n210_W_out, 
            c3_n211_W_out=> c3_n211_W_out, 
            c3_n212_W_out=> c3_n212_W_out, 
            c3_n213_W_out=> c3_n213_W_out, 
            c3_n214_W_out=> c3_n214_W_out, 
            c3_n215_W_out=> c3_n215_W_out, 
            c3_n216_W_out=> c3_n216_W_out, 
            c3_n217_W_out=> c3_n217_W_out, 
            c3_n218_W_out=> c3_n218_W_out, 
            c3_n219_W_out=> c3_n219_W_out, 
            c3_n220_W_out=> c3_n220_W_out, 
            c3_n221_W_out=> c3_n221_W_out, 
            c3_n222_W_out=> c3_n222_W_out, 
            c3_n223_W_out=> c3_n223_W_out, 
            c3_n224_W_out=> c3_n224_W_out, 
            c3_n225_W_out=> c3_n225_W_out, 
            c3_n226_W_out=> c3_n226_W_out, 
            c3_n227_W_out=> c3_n227_W_out, 
            c3_n228_W_out=> c3_n228_W_out, 
            c3_n229_W_out=> c3_n229_W_out, 
            c3_n230_W_out=> c3_n230_W_out, 
            c3_n231_W_out=> c3_n231_W_out, 
            c3_n232_W_out=> c3_n232_W_out, 
            c3_n233_W_out=> c3_n233_W_out, 
            c3_n234_W_out=> c3_n234_W_out, 
            c3_n235_W_out=> c3_n235_W_out, 
            c3_n236_W_out=> c3_n236_W_out, 
            c3_n237_W_out=> c3_n237_W_out, 
            c3_n238_W_out=> c3_n238_W_out, 
            c3_n239_W_out=> c3_n239_W_out, 
            c3_n240_W_out=> c3_n240_W_out, 
            c3_n241_W_out=> c3_n241_W_out, 
            c3_n242_W_out=> c3_n242_W_out, 
            c3_n243_W_out=> c3_n243_W_out, 
            c3_n244_W_out=> c3_n244_W_out, 
            c3_n245_W_out=> c3_n245_W_out, 
            c3_n246_W_out=> c3_n246_W_out, 
            c3_n247_W_out=> c3_n247_W_out, 
            c3_n248_W_out=> c3_n248_W_out, 
            c3_n249_W_out=> c3_n249_W_out, 
            c3_n250_W_out=> c3_n250_W_out, 
            c3_n251_W_out=> c3_n251_W_out, 
            c3_n252_W_out=> c3_n252_W_out, 
            c3_n253_W_out=> c3_n253_W_out, 
            c3_n254_W_out=> c3_n254_W_out, 
            c3_n255_W_out=> c3_n255_W_out, 
            c3_n256_W_out=> c3_n256_W_out, 
            c3_n257_W_out=> c3_n257_W_out, 
            c3_n258_W_out=> c3_n258_W_out, 
            c3_n259_W_out=> c3_n259_W_out, 
            c3_n260_W_out=> c3_n260_W_out, 
            c3_n261_W_out=> c3_n261_W_out, 
            c3_n262_W_out=> c3_n262_W_out, 
            c3_n263_W_out=> c3_n263_W_out, 
            c3_n264_W_out=> c3_n264_W_out, 
            c3_n265_W_out=> c3_n265_W_out, 
            c3_n266_W_out=> c3_n266_W_out, 
            c3_n267_W_out=> c3_n267_W_out, 
            c3_n268_W_out=> c3_n268_W_out, 
            c3_n269_W_out=> c3_n269_W_out, 
            c3_n270_W_out=> c3_n270_W_out, 
            c3_n271_W_out=> c3_n271_W_out, 
            c3_n272_W_out=> c3_n272_W_out, 
            c3_n273_W_out=> c3_n273_W_out, 
            c3_n274_W_out=> c3_n274_W_out, 
            c3_n275_W_out=> c3_n275_W_out, 
            c3_n276_W_out=> c3_n276_W_out, 
            c3_n277_W_out=> c3_n277_W_out, 
            c3_n278_W_out=> c3_n278_W_out, 
            c3_n279_W_out=> c3_n279_W_out, 
            c3_n280_W_out=> c3_n280_W_out, 
            c3_n281_W_out=> c3_n281_W_out, 
            c3_n282_W_out=> c3_n282_W_out, 
            c3_n283_W_out=> c3_n283_W_out, 
            c3_n284_W_out=> c3_n284_W_out, 
            c3_n285_W_out=> c3_n285_W_out, 
            c3_n286_W_out=> c3_n286_W_out, 
            c3_n287_W_out=> c3_n287_W_out, 
            c3_n288_W_out=> c3_n288_W_out, 
            c3_n289_W_out=> c3_n289_W_out, 
            c3_n290_W_out=> c3_n290_W_out, 
            c3_n291_W_out=> c3_n291_W_out, 
            c3_n292_W_out=> c3_n292_W_out, 
            c3_n293_W_out=> c3_n293_W_out, 
            c3_n294_W_out=> c3_n294_W_out, 
            c3_n295_W_out=> c3_n295_W_out, 
            c3_n296_W_out=> c3_n296_W_out, 
            c3_n297_W_out=> c3_n297_W_out, 
            c3_n298_W_out=> c3_n298_W_out, 
            c3_n299_W_out=> c3_n299_W_out
   );
            
camada4_inst_4: ENTITY work.camada4_Sigmoid_500neuron_8bits_300n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c4_IO_in, 
            c4_n0_W_in=> c3_n0_W_out,
            c4_n1_W_in=> c3_n1_W_out,
            c4_n2_W_in=> c3_n2_W_out,
            c4_n3_W_in=> c3_n3_W_out,
            c4_n4_W_in=> c3_n4_W_out,
            c4_n5_W_in=> c3_n5_W_out,
            c4_n6_W_in=> c3_n6_W_out,
            c4_n7_W_in=> c3_n7_W_out,
            c4_n8_W_in=> c3_n8_W_out,
            c4_n9_W_in=> c3_n9_W_out,
            c4_n10_W_in=> c3_n10_W_out,
            c4_n11_W_in=> c3_n11_W_out,
            c4_n12_W_in=> c3_n12_W_out,
            c4_n13_W_in=> c3_n13_W_out,
            c4_n14_W_in=> c3_n14_W_out,
            c4_n15_W_in=> c3_n15_W_out,
            c4_n16_W_in=> c3_n16_W_out,
            c4_n17_W_in=> c3_n17_W_out,
            c4_n18_W_in=> c3_n18_W_out,
            c4_n19_W_in=> c3_n19_W_out,
            c4_n20_W_in=> c3_n20_W_out,
            c4_n21_W_in=> c3_n21_W_out,
            c4_n22_W_in=> c3_n22_W_out,
            c4_n23_W_in=> c3_n23_W_out,
            c4_n24_W_in=> c3_n24_W_out,
            c4_n25_W_in=> c3_n25_W_out,
            c4_n26_W_in=> c3_n26_W_out,
            c4_n27_W_in=> c3_n27_W_out,
            c4_n28_W_in=> c3_n28_W_out,
            c4_n29_W_in=> c3_n29_W_out,
            c4_n30_W_in=> c3_n30_W_out,
            c4_n31_W_in=> c3_n31_W_out,
            c4_n32_W_in=> c3_n32_W_out,
            c4_n33_W_in=> c3_n33_W_out,
            c4_n34_W_in=> c3_n34_W_out,
            c4_n35_W_in=> c3_n35_W_out,
            c4_n36_W_in=> c3_n36_W_out,
            c4_n37_W_in=> c3_n37_W_out,
            c4_n38_W_in=> c3_n38_W_out,
            c4_n39_W_in=> c3_n39_W_out,
            c4_n40_W_in=> c3_n40_W_out,
            c4_n41_W_in=> c3_n41_W_out,
            c4_n42_W_in=> c3_n42_W_out,
            c4_n43_W_in=> c3_n43_W_out,
            c4_n44_W_in=> c3_n44_W_out,
            c4_n45_W_in=> c3_n45_W_out,
            c4_n46_W_in=> c3_n46_W_out,
            c4_n47_W_in=> c3_n47_W_out,
            c4_n48_W_in=> c3_n48_W_out,
            c4_n49_W_in=> c3_n49_W_out,
            c4_n50_W_in=> c3_n50_W_out,
            c4_n51_W_in=> c3_n51_W_out,
            c4_n52_W_in=> c3_n52_W_out,
            c4_n53_W_in=> c3_n53_W_out,
            c4_n54_W_in=> c3_n54_W_out,
            c4_n55_W_in=> c3_n55_W_out,
            c4_n56_W_in=> c3_n56_W_out,
            c4_n57_W_in=> c3_n57_W_out,
            c4_n58_W_in=> c3_n58_W_out,
            c4_n59_W_in=> c3_n59_W_out,
            c4_n60_W_in=> c3_n60_W_out,
            c4_n61_W_in=> c3_n61_W_out,
            c4_n62_W_in=> c3_n62_W_out,
            c4_n63_W_in=> c3_n63_W_out,
            c4_n64_W_in=> c3_n64_W_out,
            c4_n65_W_in=> c3_n65_W_out,
            c4_n66_W_in=> c3_n66_W_out,
            c4_n67_W_in=> c3_n67_W_out,
            c4_n68_W_in=> c3_n68_W_out,
            c4_n69_W_in=> c3_n69_W_out,
            c4_n70_W_in=> c3_n70_W_out,
            c4_n71_W_in=> c3_n71_W_out,
            c4_n72_W_in=> c3_n72_W_out,
            c4_n73_W_in=> c3_n73_W_out,
            c4_n74_W_in=> c3_n74_W_out,
            c4_n75_W_in=> c3_n75_W_out,
            c4_n76_W_in=> c3_n76_W_out,
            c4_n77_W_in=> c3_n77_W_out,
            c4_n78_W_in=> c3_n78_W_out,
            c4_n79_W_in=> c3_n79_W_out,
            c4_n80_W_in=> c3_n80_W_out,
            c4_n81_W_in=> c3_n81_W_out,
            c4_n82_W_in=> c3_n82_W_out,
            c4_n83_W_in=> c3_n83_W_out,
            c4_n84_W_in=> c3_n84_W_out,
            c4_n85_W_in=> c3_n85_W_out,
            c4_n86_W_in=> c3_n86_W_out,
            c4_n87_W_in=> c3_n87_W_out,
            c4_n88_W_in=> c3_n88_W_out,
            c4_n89_W_in=> c3_n89_W_out,
            c4_n90_W_in=> c3_n90_W_out,
            c4_n91_W_in=> c3_n91_W_out,
            c4_n92_W_in=> c3_n92_W_out,
            c4_n93_W_in=> c3_n93_W_out,
            c4_n94_W_in=> c3_n94_W_out,
            c4_n95_W_in=> c3_n95_W_out,
            c4_n96_W_in=> c3_n96_W_out,
            c4_n97_W_in=> c3_n97_W_out,
            c4_n98_W_in=> c3_n98_W_out,
            c4_n99_W_in=> c3_n99_W_out,
            c4_n100_W_in=> c3_n100_W_out,
            c4_n101_W_in=> c3_n101_W_out,
            c4_n102_W_in=> c3_n102_W_out,
            c4_n103_W_in=> c3_n103_W_out,
            c4_n104_W_in=> c3_n104_W_out,
            c4_n105_W_in=> c3_n105_W_out,
            c4_n106_W_in=> c3_n106_W_out,
            c4_n107_W_in=> c3_n107_W_out,
            c4_n108_W_in=> c3_n108_W_out,
            c4_n109_W_in=> c3_n109_W_out,
            c4_n110_W_in=> c3_n110_W_out,
            c4_n111_W_in=> c3_n111_W_out,
            c4_n112_W_in=> c3_n112_W_out,
            c4_n113_W_in=> c3_n113_W_out,
            c4_n114_W_in=> c3_n114_W_out,
            c4_n115_W_in=> c3_n115_W_out,
            c4_n116_W_in=> c3_n116_W_out,
            c4_n117_W_in=> c3_n117_W_out,
            c4_n118_W_in=> c3_n118_W_out,
            c4_n119_W_in=> c3_n119_W_out,
            c4_n120_W_in=> c3_n120_W_out,
            c4_n121_W_in=> c3_n121_W_out,
            c4_n122_W_in=> c3_n122_W_out,
            c4_n123_W_in=> c3_n123_W_out,
            c4_n124_W_in=> c3_n124_W_out,
            c4_n125_W_in=> c3_n125_W_out,
            c4_n126_W_in=> c3_n126_W_out,
            c4_n127_W_in=> c3_n127_W_out,
            c4_n128_W_in=> c3_n128_W_out,
            c4_n129_W_in=> c3_n129_W_out,
            c4_n130_W_in=> c3_n130_W_out,
            c4_n131_W_in=> c3_n131_W_out,
            c4_n132_W_in=> c3_n132_W_out,
            c4_n133_W_in=> c3_n133_W_out,
            c4_n134_W_in=> c3_n134_W_out,
            c4_n135_W_in=> c3_n135_W_out,
            c4_n136_W_in=> c3_n136_W_out,
            c4_n137_W_in=> c3_n137_W_out,
            c4_n138_W_in=> c3_n138_W_out,
            c4_n139_W_in=> c3_n139_W_out,
            c4_n140_W_in=> c3_n140_W_out,
            c4_n141_W_in=> c3_n141_W_out,
            c4_n142_W_in=> c3_n142_W_out,
            c4_n143_W_in=> c3_n143_W_out,
            c4_n144_W_in=> c3_n144_W_out,
            c4_n145_W_in=> c3_n145_W_out,
            c4_n146_W_in=> c3_n146_W_out,
            c4_n147_W_in=> c3_n147_W_out,
            c4_n148_W_in=> c3_n148_W_out,
            c4_n149_W_in=> c3_n149_W_out,
            c4_n150_W_in=> c3_n150_W_out,
            c4_n151_W_in=> c3_n151_W_out,
            c4_n152_W_in=> c3_n152_W_out,
            c4_n153_W_in=> c3_n153_W_out,
            c4_n154_W_in=> c3_n154_W_out,
            c4_n155_W_in=> c3_n155_W_out,
            c4_n156_W_in=> c3_n156_W_out,
            c4_n157_W_in=> c3_n157_W_out,
            c4_n158_W_in=> c3_n158_W_out,
            c4_n159_W_in=> c3_n159_W_out,
            c4_n160_W_in=> c3_n160_W_out,
            c4_n161_W_in=> c3_n161_W_out,
            c4_n162_W_in=> c3_n162_W_out,
            c4_n163_W_in=> c3_n163_W_out,
            c4_n164_W_in=> c3_n164_W_out,
            c4_n165_W_in=> c3_n165_W_out,
            c4_n166_W_in=> c3_n166_W_out,
            c4_n167_W_in=> c3_n167_W_out,
            c4_n168_W_in=> c3_n168_W_out,
            c4_n169_W_in=> c3_n169_W_out,
            c4_n170_W_in=> c3_n170_W_out,
            c4_n171_W_in=> c3_n171_W_out,
            c4_n172_W_in=> c3_n172_W_out,
            c4_n173_W_in=> c3_n173_W_out,
            c4_n174_W_in=> c3_n174_W_out,
            c4_n175_W_in=> c3_n175_W_out,
            c4_n176_W_in=> c3_n176_W_out,
            c4_n177_W_in=> c3_n177_W_out,
            c4_n178_W_in=> c3_n178_W_out,
            c4_n179_W_in=> c3_n179_W_out,
            c4_n180_W_in=> c3_n180_W_out,
            c4_n181_W_in=> c3_n181_W_out,
            c4_n182_W_in=> c3_n182_W_out,
            c4_n183_W_in=> c3_n183_W_out,
            c4_n184_W_in=> c3_n184_W_out,
            c4_n185_W_in=> c3_n185_W_out,
            c4_n186_W_in=> c3_n186_W_out,
            c4_n187_W_in=> c3_n187_W_out,
            c4_n188_W_in=> c3_n188_W_out,
            c4_n189_W_in=> c3_n189_W_out,
            c4_n190_W_in=> c3_n190_W_out,
            c4_n191_W_in=> c3_n191_W_out,
            c4_n192_W_in=> c3_n192_W_out,
            c4_n193_W_in=> c3_n193_W_out,
            c4_n194_W_in=> c3_n194_W_out,
            c4_n195_W_in=> c3_n195_W_out,
            c4_n196_W_in=> c3_n196_W_out,
            c4_n197_W_in=> c3_n197_W_out,
            c4_n198_W_in=> c3_n198_W_out,
            c4_n199_W_in=> c3_n199_W_out,
            c4_n200_W_in=> c3_n200_W_out,
            c4_n201_W_in=> c3_n201_W_out,
            c4_n202_W_in=> c3_n202_W_out,
            c4_n203_W_in=> c3_n203_W_out,
            c4_n204_W_in=> c3_n204_W_out,
            c4_n205_W_in=> c3_n205_W_out,
            c4_n206_W_in=> c3_n206_W_out,
            c4_n207_W_in=> c3_n207_W_out,
            c4_n208_W_in=> c3_n208_W_out,
            c4_n209_W_in=> c3_n209_W_out,
            c4_n210_W_in=> c3_n210_W_out,
            c4_n211_W_in=> c3_n211_W_out,
            c4_n212_W_in=> c3_n212_W_out,
            c4_n213_W_in=> c3_n213_W_out,
            c4_n214_W_in=> c3_n214_W_out,
            c4_n215_W_in=> c3_n215_W_out,
            c4_n216_W_in=> c3_n216_W_out,
            c4_n217_W_in=> c3_n217_W_out,
            c4_n218_W_in=> c3_n218_W_out,
            c4_n219_W_in=> c3_n219_W_out,
            c4_n220_W_in=> c3_n220_W_out,
            c4_n221_W_in=> c3_n221_W_out,
            c4_n222_W_in=> c3_n222_W_out,
            c4_n223_W_in=> c3_n223_W_out,
            c4_n224_W_in=> c3_n224_W_out,
            c4_n225_W_in=> c3_n225_W_out,
            c4_n226_W_in=> c3_n226_W_out,
            c4_n227_W_in=> c3_n227_W_out,
            c4_n228_W_in=> c3_n228_W_out,
            c4_n229_W_in=> c3_n229_W_out,
            c4_n230_W_in=> c3_n230_W_out,
            c4_n231_W_in=> c3_n231_W_out,
            c4_n232_W_in=> c3_n232_W_out,
            c4_n233_W_in=> c3_n233_W_out,
            c4_n234_W_in=> c3_n234_W_out,
            c4_n235_W_in=> c3_n235_W_out,
            c4_n236_W_in=> c3_n236_W_out,
            c4_n237_W_in=> c3_n237_W_out,
            c4_n238_W_in=> c3_n238_W_out,
            c4_n239_W_in=> c3_n239_W_out,
            c4_n240_W_in=> c3_n240_W_out,
            c4_n241_W_in=> c3_n241_W_out,
            c4_n242_W_in=> c3_n242_W_out,
            c4_n243_W_in=> c3_n243_W_out,
            c4_n244_W_in=> c3_n244_W_out,
            c4_n245_W_in=> c3_n245_W_out,
            c4_n246_W_in=> c3_n246_W_out,
            c4_n247_W_in=> c3_n247_W_out,
            c4_n248_W_in=> c3_n248_W_out,
            c4_n249_W_in=> c3_n249_W_out,
            c4_n250_W_in=> c3_n250_W_out,
            c4_n251_W_in=> c3_n251_W_out,
            c4_n252_W_in=> c3_n252_W_out,
            c4_n253_W_in=> c3_n253_W_out,
            c4_n254_W_in=> c3_n254_W_out,
            c4_n255_W_in=> c3_n255_W_out,
            c4_n256_W_in=> c3_n256_W_out,
            c4_n257_W_in=> c3_n257_W_out,
            c4_n258_W_in=> c3_n258_W_out,
            c4_n259_W_in=> c3_n259_W_out,
            c4_n260_W_in=> c3_n260_W_out,
            c4_n261_W_in=> c3_n261_W_out,
            c4_n262_W_in=> c3_n262_W_out,
            c4_n263_W_in=> c3_n263_W_out,
            c4_n264_W_in=> c3_n264_W_out,
            c4_n265_W_in=> c3_n265_W_out,
            c4_n266_W_in=> c3_n266_W_out,
            c4_n267_W_in=> c3_n267_W_out,
            c4_n268_W_in=> c3_n268_W_out,
            c4_n269_W_in=> c3_n269_W_out,
            c4_n270_W_in=> c3_n270_W_out,
            c4_n271_W_in=> c3_n271_W_out,
            c4_n272_W_in=> c3_n272_W_out,
            c4_n273_W_in=> c3_n273_W_out,
            c4_n274_W_in=> c3_n274_W_out,
            c4_n275_W_in=> c3_n275_W_out,
            c4_n276_W_in=> c3_n276_W_out,
            c4_n277_W_in=> c3_n277_W_out,
            c4_n278_W_in=> c3_n278_W_out,
            c4_n279_W_in=> c3_n279_W_out,
            c4_n280_W_in=> c3_n280_W_out,
            c4_n281_W_in=> c3_n281_W_out,
            c4_n282_W_in=> c3_n282_W_out,
            c4_n283_W_in=> c3_n283_W_out,
            c4_n284_W_in=> c3_n284_W_out,
            c4_n285_W_in=> c3_n285_W_out,
            c4_n286_W_in=> c3_n286_W_out,
            c4_n287_W_in=> c3_n287_W_out,
            c4_n288_W_in=> c3_n288_W_out,
            c4_n289_W_in=> c3_n289_W_out,
            c4_n290_W_in=> c3_n290_W_out,
            c4_n291_W_in=> c3_n291_W_out,
            c4_n292_W_in=> c3_n292_W_out,
            c4_n293_W_in=> c3_n293_W_out,
            c4_n294_W_in=> c3_n294_W_out,
            c4_n295_W_in=> c3_n295_W_out,
            c4_n296_W_in=> c3_n296_W_out,
            c4_n297_W_in=> c3_n297_W_out,
            c4_n298_W_in=> c3_n298_W_out,
            c4_n299_W_in=> c3_n299_W_out,
            c4_n300_W_in=> c0_n300_W_out,
            c4_n301_W_in=> c0_n301_W_out,
            c4_n302_W_in=> c0_n302_W_out,
            c4_n303_W_in=> c0_n303_W_out,
            c4_n304_W_in=> c0_n304_W_out,
            c4_n305_W_in=> c0_n305_W_out,
            c4_n306_W_in=> c0_n306_W_out,
            c4_n307_W_in=> c0_n307_W_out,
            c4_n308_W_in=> c0_n308_W_out,
            c4_n309_W_in=> c0_n309_W_out,
            c4_n310_W_in=> c0_n310_W_out,
            c4_n311_W_in=> c0_n311_W_out,
            c4_n312_W_in=> c0_n312_W_out,
            c4_n313_W_in=> c0_n313_W_out,
            c4_n314_W_in=> c0_n314_W_out,
            c4_n315_W_in=> c0_n315_W_out,
            c4_n316_W_in=> c0_n316_W_out,
            c4_n317_W_in=> c0_n317_W_out,
            c4_n318_W_in=> c0_n318_W_out,
            c4_n319_W_in=> c0_n319_W_out,
            c4_n320_W_in=> c0_n320_W_out,
            c4_n321_W_in=> c0_n321_W_out,
            c4_n322_W_in=> c0_n322_W_out,
            c4_n323_W_in=> c0_n323_W_out,
            c4_n324_W_in=> c0_n324_W_out,
            c4_n325_W_in=> c0_n325_W_out,
            c4_n326_W_in=> c0_n326_W_out,
            c4_n327_W_in=> c0_n327_W_out,
            c4_n328_W_in=> c0_n328_W_out,
            c4_n329_W_in=> c0_n329_W_out,
            c4_n330_W_in=> c0_n330_W_out,
            c4_n331_W_in=> c0_n331_W_out,
            c4_n332_W_in=> c0_n332_W_out,
            c4_n333_W_in=> c0_n333_W_out,
            c4_n334_W_in=> c0_n334_W_out,
            c4_n335_W_in=> c0_n335_W_out,
            c4_n336_W_in=> c0_n336_W_out,
            c4_n337_W_in=> c0_n337_W_out,
            c4_n338_W_in=> c0_n338_W_out,
            c4_n339_W_in=> c0_n339_W_out,
            c4_n340_W_in=> c0_n340_W_out,
            c4_n341_W_in=> c0_n341_W_out,
            c4_n342_W_in=> c0_n342_W_out,
            c4_n343_W_in=> c0_n343_W_out,
            c4_n344_W_in=> c0_n344_W_out,
            c4_n345_W_in=> c0_n345_W_out,
            c4_n346_W_in=> c0_n346_W_out,
            c4_n347_W_in=> c0_n347_W_out,
            c4_n348_W_in=> c0_n348_W_out,
            c4_n349_W_in=> c0_n349_W_out,
            c4_n350_W_in=> c0_n350_W_out,
            c4_n351_W_in=> c0_n351_W_out,
            c4_n352_W_in=> c0_n352_W_out,
            c4_n353_W_in=> c0_n353_W_out,
            c4_n354_W_in=> c0_n354_W_out,
            c4_n355_W_in=> c0_n355_W_out,
            c4_n356_W_in=> c0_n356_W_out,
            c4_n357_W_in=> c0_n357_W_out,
            c4_n358_W_in=> c0_n358_W_out,
            c4_n359_W_in=> c0_n359_W_out,
            c4_n360_W_in=> c0_n360_W_out,
            c4_n361_W_in=> c0_n361_W_out,
            c4_n362_W_in=> c0_n362_W_out,
            c4_n363_W_in=> c0_n363_W_out,
            c4_n364_W_in=> c0_n364_W_out,
            c4_n365_W_in=> c0_n365_W_out,
            c4_n366_W_in=> c0_n366_W_out,
            c4_n367_W_in=> c0_n367_W_out,
            c4_n368_W_in=> c0_n368_W_out,
            c4_n369_W_in=> c0_n369_W_out,
            c4_n370_W_in=> c0_n370_W_out,
            c4_n371_W_in=> c0_n371_W_out,
            c4_n372_W_in=> c0_n372_W_out,
            c4_n373_W_in=> c0_n373_W_out,
            c4_n374_W_in=> c0_n374_W_out,
            c4_n375_W_in=> c0_n375_W_out,
            c4_n376_W_in=> c0_n376_W_out,
            c4_n377_W_in=> c0_n377_W_out,
            c4_n378_W_in=> c0_n378_W_out,
            c4_n379_W_in=> c0_n379_W_out,
            c4_n380_W_in=> c0_n380_W_out,
            c4_n381_W_in=> c0_n381_W_out,
            c4_n382_W_in=> c0_n382_W_out,
            c4_n383_W_in=> c0_n383_W_out,
            c4_n384_W_in=> c0_n384_W_out,
            c4_n385_W_in=> c0_n385_W_out,
            c4_n386_W_in=> c0_n386_W_out,
            c4_n387_W_in=> c0_n387_W_out,
            c4_n388_W_in=> c0_n388_W_out,
            c4_n389_W_in=> c0_n389_W_out,
            c4_n390_W_in=> c0_n390_W_out,
            c4_n391_W_in=> c0_n391_W_out,
            c4_n392_W_in=> c0_n392_W_out,
            c4_n393_W_in=> c0_n393_W_out,
            c4_n394_W_in=> c0_n394_W_out,
            c4_n395_W_in=> c0_n395_W_out,
            c4_n396_W_in=> c0_n396_W_out,
            c4_n397_W_in=> c0_n397_W_out,
            c4_n398_W_in=> c0_n398_W_out,
            c4_n399_W_in=> c0_n399_W_out,
            c4_n400_W_in=> c0_n400_W_out,
            c4_n401_W_in=> c0_n401_W_out,
            c4_n402_W_in=> c0_n402_W_out,
            c4_n403_W_in=> c0_n403_W_out,
            c4_n404_W_in=> c0_n404_W_out,
            c4_n405_W_in=> c0_n405_W_out,
            c4_n406_W_in=> c0_n406_W_out,
            c4_n407_W_in=> c0_n407_W_out,
            c4_n408_W_in=> c0_n408_W_out,
            c4_n409_W_in=> c0_n409_W_out,
            c4_n410_W_in=> c0_n410_W_out,
            c4_n411_W_in=> c0_n411_W_out,
            c4_n412_W_in=> c0_n412_W_out,
            c4_n413_W_in=> c0_n413_W_out,
            c4_n414_W_in=> c0_n414_W_out,
            c4_n415_W_in=> c0_n415_W_out,
            c4_n416_W_in=> c0_n416_W_out,
            c4_n417_W_in=> c0_n417_W_out,
            c4_n418_W_in=> c0_n418_W_out,
            c4_n419_W_in=> c0_n419_W_out,
            c4_n420_W_in=> c0_n420_W_out,
            c4_n421_W_in=> c0_n421_W_out,
            c4_n422_W_in=> c0_n422_W_out,
            c4_n423_W_in=> c0_n423_W_out,
            c4_n424_W_in=> c0_n424_W_out,
            c4_n425_W_in=> c0_n425_W_out,
            c4_n426_W_in=> c0_n426_W_out,
            c4_n427_W_in=> c0_n427_W_out,
            c4_n428_W_in=> c0_n428_W_out,
            c4_n429_W_in=> c0_n429_W_out,
            c4_n430_W_in=> c0_n430_W_out,
            c4_n431_W_in=> c0_n431_W_out,
            c4_n432_W_in=> c0_n432_W_out,
            c4_n433_W_in=> c0_n433_W_out,
            c4_n434_W_in=> c0_n434_W_out,
            c4_n435_W_in=> c0_n435_W_out,
            c4_n436_W_in=> c0_n436_W_out,
            c4_n437_W_in=> c0_n437_W_out,
            c4_n438_W_in=> c0_n438_W_out,
            c4_n439_W_in=> c0_n439_W_out,
            c4_n440_W_in=> c0_n440_W_out,
            c4_n441_W_in=> c0_n441_W_out,
            c4_n442_W_in=> c0_n442_W_out,
            c4_n443_W_in=> c0_n443_W_out,
            c4_n444_W_in=> c0_n444_W_out,
            c4_n445_W_in=> c0_n445_W_out,
            c4_n446_W_in=> c0_n446_W_out,
            c4_n447_W_in=> c0_n447_W_out,
            c4_n448_W_in=> c0_n448_W_out,
            c4_n449_W_in=> c0_n449_W_out,
            c4_n450_W_in=> c0_n450_W_out,
            c4_n451_W_in=> c0_n451_W_out,
            c4_n452_W_in=> c0_n452_W_out,
            c4_n453_W_in=> c0_n453_W_out,
            c4_n454_W_in=> c0_n454_W_out,
            c4_n455_W_in=> c0_n455_W_out,
            c4_n456_W_in=> c0_n456_W_out,
            c4_n457_W_in=> c0_n457_W_out,
            c4_n458_W_in=> c0_n458_W_out,
            c4_n459_W_in=> c0_n459_W_out,
            c4_n460_W_in=> c0_n460_W_out,
            c4_n461_W_in=> c0_n461_W_out,
            c4_n462_W_in=> c0_n462_W_out,
            c4_n463_W_in=> c0_n463_W_out,
            c4_n464_W_in=> c0_n464_W_out,
            c4_n465_W_in=> c0_n465_W_out,
            c4_n466_W_in=> c0_n466_W_out,
            c4_n467_W_in=> c0_n467_W_out,
            c4_n468_W_in=> c0_n468_W_out,
            c4_n469_W_in=> c0_n469_W_out,
            c4_n470_W_in=> c0_n470_W_out,
            c4_n471_W_in=> c0_n471_W_out,
            c4_n472_W_in=> c0_n472_W_out,
            c4_n473_W_in=> c0_n473_W_out,
            c4_n474_W_in=> c0_n474_W_out,
            c4_n475_W_in=> c0_n475_W_out,
            c4_n476_W_in=> c0_n476_W_out,
            c4_n477_W_in=> c0_n477_W_out,
            c4_n478_W_in=> c0_n478_W_out,
            c4_n479_W_in=> c0_n479_W_out,
            c4_n480_W_in=> c0_n480_W_out,
            c4_n481_W_in=> c0_n481_W_out,
            c4_n482_W_in=> c0_n482_W_out,
            c4_n483_W_in=> c0_n483_W_out,
            c4_n484_W_in=> c0_n484_W_out,
            c4_n485_W_in=> c0_n485_W_out,
            c4_n486_W_in=> c0_n486_W_out,
            c4_n487_W_in=> c0_n487_W_out,
            c4_n488_W_in=> c0_n488_W_out,
            c4_n489_W_in=> c0_n489_W_out,
            c4_n490_W_in=> c0_n490_W_out,
            c4_n491_W_in=> c0_n491_W_out,
            c4_n492_W_in=> c0_n492_W_out,
            c4_n493_W_in=> c0_n493_W_out,
            c4_n494_W_in=> c0_n494_W_out,
            c4_n495_W_in=> c0_n495_W_out,
            c4_n496_W_in=> c0_n496_W_out,
            c4_n497_W_in=> c0_n497_W_out,
            c4_n498_W_in=> c0_n498_W_out,
            c4_n499_W_in=> c0_n499_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c4_n0_IO_out=> c4_n0_IO_out, 
            c4_n1_IO_out=> c4_n1_IO_out, 
            c4_n2_IO_out=> c4_n2_IO_out, 
            c4_n3_IO_out=> c4_n3_IO_out, 
            c4_n4_IO_out=> c4_n4_IO_out, 
            c4_n5_IO_out=> c4_n5_IO_out, 
            c4_n6_IO_out=> c4_n6_IO_out, 
            c4_n7_IO_out=> c4_n7_IO_out, 
            c4_n8_IO_out=> c4_n8_IO_out, 
            c4_n9_IO_out=> c4_n9_IO_out, 
            c4_n10_IO_out=> c4_n10_IO_out, 
            c4_n11_IO_out=> c4_n11_IO_out, 
            c4_n12_IO_out=> c4_n12_IO_out, 
            c4_n13_IO_out=> c4_n13_IO_out, 
            c4_n14_IO_out=> c4_n14_IO_out, 
            c4_n15_IO_out=> c4_n15_IO_out, 
            c4_n16_IO_out=> c4_n16_IO_out, 
            c4_n17_IO_out=> c4_n17_IO_out, 
            c4_n18_IO_out=> c4_n18_IO_out, 
            c4_n19_IO_out=> c4_n19_IO_out, 
            c4_n20_IO_out=> c4_n20_IO_out, 
            c4_n21_IO_out=> c4_n21_IO_out, 
            c4_n22_IO_out=> c4_n22_IO_out, 
            c4_n23_IO_out=> c4_n23_IO_out, 
            c4_n24_IO_out=> c4_n24_IO_out, 
            c4_n25_IO_out=> c4_n25_IO_out, 
            c4_n26_IO_out=> c4_n26_IO_out, 
            c4_n27_IO_out=> c4_n27_IO_out, 
            c4_n28_IO_out=> c4_n28_IO_out, 
            c4_n29_IO_out=> c4_n29_IO_out, 
            c4_n30_IO_out=> c4_n30_IO_out, 
            c4_n31_IO_out=> c4_n31_IO_out, 
            c4_n32_IO_out=> c4_n32_IO_out, 
            c4_n33_IO_out=> c4_n33_IO_out, 
            c4_n34_IO_out=> c4_n34_IO_out, 
            c4_n35_IO_out=> c4_n35_IO_out, 
            c4_n36_IO_out=> c4_n36_IO_out, 
            c4_n37_IO_out=> c4_n37_IO_out, 
            c4_n38_IO_out=> c4_n38_IO_out, 
            c4_n39_IO_out=> c4_n39_IO_out, 
            c4_n40_IO_out=> c4_n40_IO_out, 
            c4_n41_IO_out=> c4_n41_IO_out, 
            c4_n42_IO_out=> c4_n42_IO_out, 
            c4_n43_IO_out=> c4_n43_IO_out, 
            c4_n44_IO_out=> c4_n44_IO_out, 
            c4_n45_IO_out=> c4_n45_IO_out, 
            c4_n46_IO_out=> c4_n46_IO_out, 
            c4_n47_IO_out=> c4_n47_IO_out, 
            c4_n48_IO_out=> c4_n48_IO_out, 
            c4_n49_IO_out=> c4_n49_IO_out, 
            c4_n50_IO_out=> c4_n50_IO_out, 
            c4_n51_IO_out=> c4_n51_IO_out, 
            c4_n52_IO_out=> c4_n52_IO_out, 
            c4_n53_IO_out=> c4_n53_IO_out, 
            c4_n54_IO_out=> c4_n54_IO_out, 
            c4_n55_IO_out=> c4_n55_IO_out, 
            c4_n56_IO_out=> c4_n56_IO_out, 
            c4_n57_IO_out=> c4_n57_IO_out, 
            c4_n58_IO_out=> c4_n58_IO_out, 
            c4_n59_IO_out=> c4_n59_IO_out, 
            c4_n60_IO_out=> c4_n60_IO_out, 
            c4_n61_IO_out=> c4_n61_IO_out, 
            c4_n62_IO_out=> c4_n62_IO_out, 
            c4_n63_IO_out=> c4_n63_IO_out, 
            c4_n64_IO_out=> c4_n64_IO_out, 
            c4_n65_IO_out=> c4_n65_IO_out, 
            c4_n66_IO_out=> c4_n66_IO_out, 
            c4_n67_IO_out=> c4_n67_IO_out, 
            c4_n68_IO_out=> c4_n68_IO_out, 
            c4_n69_IO_out=> c4_n69_IO_out, 
            c4_n70_IO_out=> c4_n70_IO_out, 
            c4_n71_IO_out=> c4_n71_IO_out, 
            c4_n72_IO_out=> c4_n72_IO_out, 
            c4_n73_IO_out=> c4_n73_IO_out, 
            c4_n74_IO_out=> c4_n74_IO_out, 
            c4_n75_IO_out=> c4_n75_IO_out, 
            c4_n76_IO_out=> c4_n76_IO_out, 
            c4_n77_IO_out=> c4_n77_IO_out, 
            c4_n78_IO_out=> c4_n78_IO_out, 
            c4_n79_IO_out=> c4_n79_IO_out, 
            c4_n80_IO_out=> c4_n80_IO_out, 
            c4_n81_IO_out=> c4_n81_IO_out, 
            c4_n82_IO_out=> c4_n82_IO_out, 
            c4_n83_IO_out=> c4_n83_IO_out, 
            c4_n84_IO_out=> c4_n84_IO_out, 
            c4_n85_IO_out=> c4_n85_IO_out, 
            c4_n86_IO_out=> c4_n86_IO_out, 
            c4_n87_IO_out=> c4_n87_IO_out, 
            c4_n88_IO_out=> c4_n88_IO_out, 
            c4_n89_IO_out=> c4_n89_IO_out, 
            c4_n90_IO_out=> c4_n90_IO_out, 
            c4_n91_IO_out=> c4_n91_IO_out, 
            c4_n92_IO_out=> c4_n92_IO_out, 
            c4_n93_IO_out=> c4_n93_IO_out, 
            c4_n94_IO_out=> c4_n94_IO_out, 
            c4_n95_IO_out=> c4_n95_IO_out, 
            c4_n96_IO_out=> c4_n96_IO_out, 
            c4_n97_IO_out=> c4_n97_IO_out, 
            c4_n98_IO_out=> c4_n98_IO_out, 
            c4_n99_IO_out=> c4_n99_IO_out, 
            c4_n100_IO_out=> c4_n100_IO_out, 
            c4_n101_IO_out=> c4_n101_IO_out, 
            c4_n102_IO_out=> c4_n102_IO_out, 
            c4_n103_IO_out=> c4_n103_IO_out, 
            c4_n104_IO_out=> c4_n104_IO_out, 
            c4_n105_IO_out=> c4_n105_IO_out, 
            c4_n106_IO_out=> c4_n106_IO_out, 
            c4_n107_IO_out=> c4_n107_IO_out, 
            c4_n108_IO_out=> c4_n108_IO_out, 
            c4_n109_IO_out=> c4_n109_IO_out, 
            c4_n110_IO_out=> c4_n110_IO_out, 
            c4_n111_IO_out=> c4_n111_IO_out, 
            c4_n112_IO_out=> c4_n112_IO_out, 
            c4_n113_IO_out=> c4_n113_IO_out, 
            c4_n114_IO_out=> c4_n114_IO_out, 
            c4_n115_IO_out=> c4_n115_IO_out, 
            c4_n116_IO_out=> c4_n116_IO_out, 
            c4_n117_IO_out=> c4_n117_IO_out, 
            c4_n118_IO_out=> c4_n118_IO_out, 
            c4_n119_IO_out=> c4_n119_IO_out, 
            c4_n120_IO_out=> c4_n120_IO_out, 
            c4_n121_IO_out=> c4_n121_IO_out, 
            c4_n122_IO_out=> c4_n122_IO_out, 
            c4_n123_IO_out=> c4_n123_IO_out, 
            c4_n124_IO_out=> c4_n124_IO_out, 
            c4_n125_IO_out=> c4_n125_IO_out, 
            c4_n126_IO_out=> c4_n126_IO_out, 
            c4_n127_IO_out=> c4_n127_IO_out, 
            c4_n128_IO_out=> c4_n128_IO_out, 
            c4_n129_IO_out=> c4_n129_IO_out, 
            c4_n130_IO_out=> c4_n130_IO_out, 
            c4_n131_IO_out=> c4_n131_IO_out, 
            c4_n132_IO_out=> c4_n132_IO_out, 
            c4_n133_IO_out=> c4_n133_IO_out, 
            c4_n134_IO_out=> c4_n134_IO_out, 
            c4_n135_IO_out=> c4_n135_IO_out, 
            c4_n136_IO_out=> c4_n136_IO_out, 
            c4_n137_IO_out=> c4_n137_IO_out, 
            c4_n138_IO_out=> c4_n138_IO_out, 
            c4_n139_IO_out=> c4_n139_IO_out, 
            c4_n140_IO_out=> c4_n140_IO_out, 
            c4_n141_IO_out=> c4_n141_IO_out, 
            c4_n142_IO_out=> c4_n142_IO_out, 
            c4_n143_IO_out=> c4_n143_IO_out, 
            c4_n144_IO_out=> c4_n144_IO_out, 
            c4_n145_IO_out=> c4_n145_IO_out, 
            c4_n146_IO_out=> c4_n146_IO_out, 
            c4_n147_IO_out=> c4_n147_IO_out, 
            c4_n148_IO_out=> c4_n148_IO_out, 
            c4_n149_IO_out=> c4_n149_IO_out, 
            c4_n150_IO_out=> c4_n150_IO_out, 
            c4_n151_IO_out=> c4_n151_IO_out, 
            c4_n152_IO_out=> c4_n152_IO_out, 
            c4_n153_IO_out=> c4_n153_IO_out, 
            c4_n154_IO_out=> c4_n154_IO_out, 
            c4_n155_IO_out=> c4_n155_IO_out, 
            c4_n156_IO_out=> c4_n156_IO_out, 
            c4_n157_IO_out=> c4_n157_IO_out, 
            c4_n158_IO_out=> c4_n158_IO_out, 
            c4_n159_IO_out=> c4_n159_IO_out, 
            c4_n160_IO_out=> c4_n160_IO_out, 
            c4_n161_IO_out=> c4_n161_IO_out, 
            c4_n162_IO_out=> c4_n162_IO_out, 
            c4_n163_IO_out=> c4_n163_IO_out, 
            c4_n164_IO_out=> c4_n164_IO_out, 
            c4_n165_IO_out=> c4_n165_IO_out, 
            c4_n166_IO_out=> c4_n166_IO_out, 
            c4_n167_IO_out=> c4_n167_IO_out, 
            c4_n168_IO_out=> c4_n168_IO_out, 
            c4_n169_IO_out=> c4_n169_IO_out, 
            c4_n170_IO_out=> c4_n170_IO_out, 
            c4_n171_IO_out=> c4_n171_IO_out, 
            c4_n172_IO_out=> c4_n172_IO_out, 
            c4_n173_IO_out=> c4_n173_IO_out, 
            c4_n174_IO_out=> c4_n174_IO_out, 
            c4_n175_IO_out=> c4_n175_IO_out, 
            c4_n176_IO_out=> c4_n176_IO_out, 
            c4_n177_IO_out=> c4_n177_IO_out, 
            c4_n178_IO_out=> c4_n178_IO_out, 
            c4_n179_IO_out=> c4_n179_IO_out, 
            c4_n180_IO_out=> c4_n180_IO_out, 
            c4_n181_IO_out=> c4_n181_IO_out, 
            c4_n182_IO_out=> c4_n182_IO_out, 
            c4_n183_IO_out=> c4_n183_IO_out, 
            c4_n184_IO_out=> c4_n184_IO_out, 
            c4_n185_IO_out=> c4_n185_IO_out, 
            c4_n186_IO_out=> c4_n186_IO_out, 
            c4_n187_IO_out=> c4_n187_IO_out, 
            c4_n188_IO_out=> c4_n188_IO_out, 
            c4_n189_IO_out=> c4_n189_IO_out, 
            c4_n190_IO_out=> c4_n190_IO_out, 
            c4_n191_IO_out=> c4_n191_IO_out, 
            c4_n192_IO_out=> c4_n192_IO_out, 
            c4_n193_IO_out=> c4_n193_IO_out, 
            c4_n194_IO_out=> c4_n194_IO_out, 
            c4_n195_IO_out=> c4_n195_IO_out, 
            c4_n196_IO_out=> c4_n196_IO_out, 
            c4_n197_IO_out=> c4_n197_IO_out, 
            c4_n198_IO_out=> c4_n198_IO_out, 
            c4_n199_IO_out=> c4_n199_IO_out, 
            c4_n200_IO_out=> c4_n200_IO_out, 
            c4_n201_IO_out=> c4_n201_IO_out, 
            c4_n202_IO_out=> c4_n202_IO_out, 
            c4_n203_IO_out=> c4_n203_IO_out, 
            c4_n204_IO_out=> c4_n204_IO_out, 
            c4_n205_IO_out=> c4_n205_IO_out, 
            c4_n206_IO_out=> c4_n206_IO_out, 
            c4_n207_IO_out=> c4_n207_IO_out, 
            c4_n208_IO_out=> c4_n208_IO_out, 
            c4_n209_IO_out=> c4_n209_IO_out, 
            c4_n210_IO_out=> c4_n210_IO_out, 
            c4_n211_IO_out=> c4_n211_IO_out, 
            c4_n212_IO_out=> c4_n212_IO_out, 
            c4_n213_IO_out=> c4_n213_IO_out, 
            c4_n214_IO_out=> c4_n214_IO_out, 
            c4_n215_IO_out=> c4_n215_IO_out, 
            c4_n216_IO_out=> c4_n216_IO_out, 
            c4_n217_IO_out=> c4_n217_IO_out, 
            c4_n218_IO_out=> c4_n218_IO_out, 
            c4_n219_IO_out=> c4_n219_IO_out, 
            c4_n220_IO_out=> c4_n220_IO_out, 
            c4_n221_IO_out=> c4_n221_IO_out, 
            c4_n222_IO_out=> c4_n222_IO_out, 
            c4_n223_IO_out=> c4_n223_IO_out, 
            c4_n224_IO_out=> c4_n224_IO_out, 
            c4_n225_IO_out=> c4_n225_IO_out, 
            c4_n226_IO_out=> c4_n226_IO_out, 
            c4_n227_IO_out=> c4_n227_IO_out, 
            c4_n228_IO_out=> c4_n228_IO_out, 
            c4_n229_IO_out=> c4_n229_IO_out, 
            c4_n230_IO_out=> c4_n230_IO_out, 
            c4_n231_IO_out=> c4_n231_IO_out, 
            c4_n232_IO_out=> c4_n232_IO_out, 
            c4_n233_IO_out=> c4_n233_IO_out, 
            c4_n234_IO_out=> c4_n234_IO_out, 
            c4_n235_IO_out=> c4_n235_IO_out, 
            c4_n236_IO_out=> c4_n236_IO_out, 
            c4_n237_IO_out=> c4_n237_IO_out, 
            c4_n238_IO_out=> c4_n238_IO_out, 
            c4_n239_IO_out=> c4_n239_IO_out, 
            c4_n240_IO_out=> c4_n240_IO_out, 
            c4_n241_IO_out=> c4_n241_IO_out, 
            c4_n242_IO_out=> c4_n242_IO_out, 
            c4_n243_IO_out=> c4_n243_IO_out, 
            c4_n244_IO_out=> c4_n244_IO_out, 
            c4_n245_IO_out=> c4_n245_IO_out, 
            c4_n246_IO_out=> c4_n246_IO_out, 
            c4_n247_IO_out=> c4_n247_IO_out, 
            c4_n248_IO_out=> c4_n248_IO_out, 
            c4_n249_IO_out=> c4_n249_IO_out, 
            c4_n250_IO_out=> c4_n250_IO_out, 
            c4_n251_IO_out=> c4_n251_IO_out, 
            c4_n252_IO_out=> c4_n252_IO_out, 
            c4_n253_IO_out=> c4_n253_IO_out, 
            c4_n254_IO_out=> c4_n254_IO_out, 
            c4_n255_IO_out=> c4_n255_IO_out, 
            c4_n256_IO_out=> c4_n256_IO_out, 
            c4_n257_IO_out=> c4_n257_IO_out, 
            c4_n258_IO_out=> c4_n258_IO_out, 
            c4_n259_IO_out=> c4_n259_IO_out, 
            c4_n260_IO_out=> c4_n260_IO_out, 
            c4_n261_IO_out=> c4_n261_IO_out, 
            c4_n262_IO_out=> c4_n262_IO_out, 
            c4_n263_IO_out=> c4_n263_IO_out, 
            c4_n264_IO_out=> c4_n264_IO_out, 
            c4_n265_IO_out=> c4_n265_IO_out, 
            c4_n266_IO_out=> c4_n266_IO_out, 
            c4_n267_IO_out=> c4_n267_IO_out, 
            c4_n268_IO_out=> c4_n268_IO_out, 
            c4_n269_IO_out=> c4_n269_IO_out, 
            c4_n270_IO_out=> c4_n270_IO_out, 
            c4_n271_IO_out=> c4_n271_IO_out, 
            c4_n272_IO_out=> c4_n272_IO_out, 
            c4_n273_IO_out=> c4_n273_IO_out, 
            c4_n274_IO_out=> c4_n274_IO_out, 
            c4_n275_IO_out=> c4_n275_IO_out, 
            c4_n276_IO_out=> c4_n276_IO_out, 
            c4_n277_IO_out=> c4_n277_IO_out, 
            c4_n278_IO_out=> c4_n278_IO_out, 
            c4_n279_IO_out=> c4_n279_IO_out, 
            c4_n280_IO_out=> c4_n280_IO_out, 
            c4_n281_IO_out=> c4_n281_IO_out, 
            c4_n282_IO_out=> c4_n282_IO_out, 
            c4_n283_IO_out=> c4_n283_IO_out, 
            c4_n284_IO_out=> c4_n284_IO_out, 
            c4_n285_IO_out=> c4_n285_IO_out, 
            c4_n286_IO_out=> c4_n286_IO_out, 
            c4_n287_IO_out=> c4_n287_IO_out, 
            c4_n288_IO_out=> c4_n288_IO_out, 
            c4_n289_IO_out=> c4_n289_IO_out, 
            c4_n290_IO_out=> c4_n290_IO_out, 
            c4_n291_IO_out=> c4_n291_IO_out, 
            c4_n292_IO_out=> c4_n292_IO_out, 
            c4_n293_IO_out=> c4_n293_IO_out, 
            c4_n294_IO_out=> c4_n294_IO_out, 
            c4_n295_IO_out=> c4_n295_IO_out, 
            c4_n296_IO_out=> c4_n296_IO_out, 
            c4_n297_IO_out=> c4_n297_IO_out, 
            c4_n298_IO_out=> c4_n298_IO_out, 
            c4_n299_IO_out=> c4_n299_IO_out, 
            c4_n300_IO_out=> c4_n300_IO_out, 
            c4_n301_IO_out=> c4_n301_IO_out, 
            c4_n302_IO_out=> c4_n302_IO_out, 
            c4_n303_IO_out=> c4_n303_IO_out, 
            c4_n304_IO_out=> c4_n304_IO_out, 
            c4_n305_IO_out=> c4_n305_IO_out, 
            c4_n306_IO_out=> c4_n306_IO_out, 
            c4_n307_IO_out=> c4_n307_IO_out, 
            c4_n308_IO_out=> c4_n308_IO_out, 
            c4_n309_IO_out=> c4_n309_IO_out, 
            c4_n310_IO_out=> c4_n310_IO_out, 
            c4_n311_IO_out=> c4_n311_IO_out, 
            c4_n312_IO_out=> c4_n312_IO_out, 
            c4_n313_IO_out=> c4_n313_IO_out, 
            c4_n314_IO_out=> c4_n314_IO_out, 
            c4_n315_IO_out=> c4_n315_IO_out, 
            c4_n316_IO_out=> c4_n316_IO_out, 
            c4_n317_IO_out=> c4_n317_IO_out, 
            c4_n318_IO_out=> c4_n318_IO_out, 
            c4_n319_IO_out=> c4_n319_IO_out, 
            c4_n320_IO_out=> c4_n320_IO_out, 
            c4_n321_IO_out=> c4_n321_IO_out, 
            c4_n322_IO_out=> c4_n322_IO_out, 
            c4_n323_IO_out=> c4_n323_IO_out, 
            c4_n324_IO_out=> c4_n324_IO_out, 
            c4_n325_IO_out=> c4_n325_IO_out, 
            c4_n326_IO_out=> c4_n326_IO_out, 
            c4_n327_IO_out=> c4_n327_IO_out, 
            c4_n328_IO_out=> c4_n328_IO_out, 
            c4_n329_IO_out=> c4_n329_IO_out, 
            c4_n330_IO_out=> c4_n330_IO_out, 
            c4_n331_IO_out=> c4_n331_IO_out, 
            c4_n332_IO_out=> c4_n332_IO_out, 
            c4_n333_IO_out=> c4_n333_IO_out, 
            c4_n334_IO_out=> c4_n334_IO_out, 
            c4_n335_IO_out=> c4_n335_IO_out, 
            c4_n336_IO_out=> c4_n336_IO_out, 
            c4_n337_IO_out=> c4_n337_IO_out, 
            c4_n338_IO_out=> c4_n338_IO_out, 
            c4_n339_IO_out=> c4_n339_IO_out, 
            c4_n340_IO_out=> c4_n340_IO_out, 
            c4_n341_IO_out=> c4_n341_IO_out, 
            c4_n342_IO_out=> c4_n342_IO_out, 
            c4_n343_IO_out=> c4_n343_IO_out, 
            c4_n344_IO_out=> c4_n344_IO_out, 
            c4_n345_IO_out=> c4_n345_IO_out, 
            c4_n346_IO_out=> c4_n346_IO_out, 
            c4_n347_IO_out=> c4_n347_IO_out, 
            c4_n348_IO_out=> c4_n348_IO_out, 
            c4_n349_IO_out=> c4_n349_IO_out, 
            c4_n350_IO_out=> c4_n350_IO_out, 
            c4_n351_IO_out=> c4_n351_IO_out, 
            c4_n352_IO_out=> c4_n352_IO_out, 
            c4_n353_IO_out=> c4_n353_IO_out, 
            c4_n354_IO_out=> c4_n354_IO_out, 
            c4_n355_IO_out=> c4_n355_IO_out, 
            c4_n356_IO_out=> c4_n356_IO_out, 
            c4_n357_IO_out=> c4_n357_IO_out, 
            c4_n358_IO_out=> c4_n358_IO_out, 
            c4_n359_IO_out=> c4_n359_IO_out, 
            c4_n360_IO_out=> c4_n360_IO_out, 
            c4_n361_IO_out=> c4_n361_IO_out, 
            c4_n362_IO_out=> c4_n362_IO_out, 
            c4_n363_IO_out=> c4_n363_IO_out, 
            c4_n364_IO_out=> c4_n364_IO_out, 
            c4_n365_IO_out=> c4_n365_IO_out, 
            c4_n366_IO_out=> c4_n366_IO_out, 
            c4_n367_IO_out=> c4_n367_IO_out, 
            c4_n368_IO_out=> c4_n368_IO_out, 
            c4_n369_IO_out=> c4_n369_IO_out, 
            c4_n370_IO_out=> c4_n370_IO_out, 
            c4_n371_IO_out=> c4_n371_IO_out, 
            c4_n372_IO_out=> c4_n372_IO_out, 
            c4_n373_IO_out=> c4_n373_IO_out, 
            c4_n374_IO_out=> c4_n374_IO_out, 
            c4_n375_IO_out=> c4_n375_IO_out, 
            c4_n376_IO_out=> c4_n376_IO_out, 
            c4_n377_IO_out=> c4_n377_IO_out, 
            c4_n378_IO_out=> c4_n378_IO_out, 
            c4_n379_IO_out=> c4_n379_IO_out, 
            c4_n380_IO_out=> c4_n380_IO_out, 
            c4_n381_IO_out=> c4_n381_IO_out, 
            c4_n382_IO_out=> c4_n382_IO_out, 
            c4_n383_IO_out=> c4_n383_IO_out, 
            c4_n384_IO_out=> c4_n384_IO_out, 
            c4_n385_IO_out=> c4_n385_IO_out, 
            c4_n386_IO_out=> c4_n386_IO_out, 
            c4_n387_IO_out=> c4_n387_IO_out, 
            c4_n388_IO_out=> c4_n388_IO_out, 
            c4_n389_IO_out=> c4_n389_IO_out, 
            c4_n390_IO_out=> c4_n390_IO_out, 
            c4_n391_IO_out=> c4_n391_IO_out, 
            c4_n392_IO_out=> c4_n392_IO_out, 
            c4_n393_IO_out=> c4_n393_IO_out, 
            c4_n394_IO_out=> c4_n394_IO_out, 
            c4_n395_IO_out=> c4_n395_IO_out, 
            c4_n396_IO_out=> c4_n396_IO_out, 
            c4_n397_IO_out=> c4_n397_IO_out, 
            c4_n398_IO_out=> c4_n398_IO_out, 
            c4_n399_IO_out=> c4_n399_IO_out, 
            c4_n400_IO_out=> c4_n400_IO_out, 
            c4_n401_IO_out=> c4_n401_IO_out, 
            c4_n402_IO_out=> c4_n402_IO_out, 
            c4_n403_IO_out=> c4_n403_IO_out, 
            c4_n404_IO_out=> c4_n404_IO_out, 
            c4_n405_IO_out=> c4_n405_IO_out, 
            c4_n406_IO_out=> c4_n406_IO_out, 
            c4_n407_IO_out=> c4_n407_IO_out, 
            c4_n408_IO_out=> c4_n408_IO_out, 
            c4_n409_IO_out=> c4_n409_IO_out, 
            c4_n410_IO_out=> c4_n410_IO_out, 
            c4_n411_IO_out=> c4_n411_IO_out, 
            c4_n412_IO_out=> c4_n412_IO_out, 
            c4_n413_IO_out=> c4_n413_IO_out, 
            c4_n414_IO_out=> c4_n414_IO_out, 
            c4_n415_IO_out=> c4_n415_IO_out, 
            c4_n416_IO_out=> c4_n416_IO_out, 
            c4_n417_IO_out=> c4_n417_IO_out, 
            c4_n418_IO_out=> c4_n418_IO_out, 
            c4_n419_IO_out=> c4_n419_IO_out, 
            c4_n420_IO_out=> c4_n420_IO_out, 
            c4_n421_IO_out=> c4_n421_IO_out, 
            c4_n422_IO_out=> c4_n422_IO_out, 
            c4_n423_IO_out=> c4_n423_IO_out, 
            c4_n424_IO_out=> c4_n424_IO_out, 
            c4_n425_IO_out=> c4_n425_IO_out, 
            c4_n426_IO_out=> c4_n426_IO_out, 
            c4_n427_IO_out=> c4_n427_IO_out, 
            c4_n428_IO_out=> c4_n428_IO_out, 
            c4_n429_IO_out=> c4_n429_IO_out, 
            c4_n430_IO_out=> c4_n430_IO_out, 
            c4_n431_IO_out=> c4_n431_IO_out, 
            c4_n432_IO_out=> c4_n432_IO_out, 
            c4_n433_IO_out=> c4_n433_IO_out, 
            c4_n434_IO_out=> c4_n434_IO_out, 
            c4_n435_IO_out=> c4_n435_IO_out, 
            c4_n436_IO_out=> c4_n436_IO_out, 
            c4_n437_IO_out=> c4_n437_IO_out, 
            c4_n438_IO_out=> c4_n438_IO_out, 
            c4_n439_IO_out=> c4_n439_IO_out, 
            c4_n440_IO_out=> c4_n440_IO_out, 
            c4_n441_IO_out=> c4_n441_IO_out, 
            c4_n442_IO_out=> c4_n442_IO_out, 
            c4_n443_IO_out=> c4_n443_IO_out, 
            c4_n444_IO_out=> c4_n444_IO_out, 
            c4_n445_IO_out=> c4_n445_IO_out, 
            c4_n446_IO_out=> c4_n446_IO_out, 
            c4_n447_IO_out=> c4_n447_IO_out, 
            c4_n448_IO_out=> c4_n448_IO_out, 
            c4_n449_IO_out=> c4_n449_IO_out, 
            c4_n450_IO_out=> c4_n450_IO_out, 
            c4_n451_IO_out=> c4_n451_IO_out, 
            c4_n452_IO_out=> c4_n452_IO_out, 
            c4_n453_IO_out=> c4_n453_IO_out, 
            c4_n454_IO_out=> c4_n454_IO_out, 
            c4_n455_IO_out=> c4_n455_IO_out, 
            c4_n456_IO_out=> c4_n456_IO_out, 
            c4_n457_IO_out=> c4_n457_IO_out, 
            c4_n458_IO_out=> c4_n458_IO_out, 
            c4_n459_IO_out=> c4_n459_IO_out, 
            c4_n460_IO_out=> c4_n460_IO_out, 
            c4_n461_IO_out=> c4_n461_IO_out, 
            c4_n462_IO_out=> c4_n462_IO_out, 
            c4_n463_IO_out=> c4_n463_IO_out, 
            c4_n464_IO_out=> c4_n464_IO_out, 
            c4_n465_IO_out=> c4_n465_IO_out, 
            c4_n466_IO_out=> c4_n466_IO_out, 
            c4_n467_IO_out=> c4_n467_IO_out, 
            c4_n468_IO_out=> c4_n468_IO_out, 
            c4_n469_IO_out=> c4_n469_IO_out, 
            c4_n470_IO_out=> c4_n470_IO_out, 
            c4_n471_IO_out=> c4_n471_IO_out, 
            c4_n472_IO_out=> c4_n472_IO_out, 
            c4_n473_IO_out=> c4_n473_IO_out, 
            c4_n474_IO_out=> c4_n474_IO_out, 
            c4_n475_IO_out=> c4_n475_IO_out, 
            c4_n476_IO_out=> c4_n476_IO_out, 
            c4_n477_IO_out=> c4_n477_IO_out, 
            c4_n478_IO_out=> c4_n478_IO_out, 
            c4_n479_IO_out=> c4_n479_IO_out, 
            c4_n480_IO_out=> c4_n480_IO_out, 
            c4_n481_IO_out=> c4_n481_IO_out, 
            c4_n482_IO_out=> c4_n482_IO_out, 
            c4_n483_IO_out=> c4_n483_IO_out, 
            c4_n484_IO_out=> c4_n484_IO_out, 
            c4_n485_IO_out=> c4_n485_IO_out, 
            c4_n486_IO_out=> c4_n486_IO_out, 
            c4_n487_IO_out=> c4_n487_IO_out, 
            c4_n488_IO_out=> c4_n488_IO_out, 
            c4_n489_IO_out=> c4_n489_IO_out, 
            c4_n490_IO_out=> c4_n490_IO_out, 
            c4_n491_IO_out=> c4_n491_IO_out, 
            c4_n492_IO_out=> c4_n492_IO_out, 
            c4_n493_IO_out=> c4_n493_IO_out, 
            c4_n494_IO_out=> c4_n494_IO_out, 
            c4_n495_IO_out=> c4_n495_IO_out, 
            c4_n496_IO_out=> c4_n496_IO_out, 
            c4_n497_IO_out=> c4_n497_IO_out, 
            c4_n498_IO_out=> c4_n498_IO_out, 
            c4_n499_IO_out=> c4_n499_IO_out
   );
            
END ARCHITECTURE;
