LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada1_ReLU_50neuron_8bits_100n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c1_n0_bias, c1_n1_bias, c1_n2_bias, c1_n3_bias, c1_n4_bias, c1_n5_bias, c1_n6_bias, c1_n7_bias, c1_n8_bias, c1_n9_bias, c1_n10_bias, c1_n11_bias, c1_n12_bias, c1_n13_bias, c1_n14_bias, c1_n15_bias, c1_n16_bias, c1_n17_bias, c1_n18_bias, c1_n19_bias, c1_n20_bias, c1_n21_bias, c1_n22_bias, c1_n23_bias, c1_n24_bias, c1_n25_bias, c1_n26_bias, c1_n27_bias, c1_n28_bias, c1_n29_bias, c1_n30_bias, c1_n31_bias, c1_n32_bias, c1_n33_bias, c1_n34_bias, c1_n35_bias, c1_n36_bias, c1_n37_bias, c1_n38_bias, c1_n39_bias, c1_n40_bias, c1_n41_bias, c1_n42_bias, c1_n43_bias, c1_n44_bias, c1_n45_bias, c1_n46_bias, c1_n47_bias, c1_n48_bias, c1_n49_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, c1_n0_w1, c1_n0_w2, c1_n0_w3, c1_n0_w4, c1_n0_w5, c1_n0_w6, c1_n0_w7, c1_n0_w8, c1_n0_w9, c1_n0_w10, c1_n0_w11, c1_n0_w12, c1_n0_w13, c1_n0_w14, c1_n0_w15, c1_n0_w16, c1_n0_w17, c1_n0_w18, c1_n0_w19, c1_n0_w20, c1_n0_w21, c1_n0_w22, c1_n0_w23, c1_n0_w24, c1_n0_w25, c1_n0_w26, c1_n0_w27, c1_n0_w28, c1_n0_w29, c1_n0_w30, c1_n0_w31, c1_n0_w32, c1_n0_w33, c1_n0_w34, c1_n0_w35, c1_n0_w36, c1_n0_w37, c1_n0_w38, c1_n0_w39, c1_n0_w40, c1_n0_w41, c1_n0_w42, c1_n0_w43, c1_n0_w44, c1_n0_w45, c1_n0_w46, c1_n0_w47, c1_n0_w48, c1_n0_w49, c1_n0_w50, c1_n0_w51, c1_n0_w52, c1_n0_w53, c1_n0_w54, c1_n0_w55, c1_n0_w56, c1_n0_w57, c1_n0_w58, c1_n0_w59, c1_n0_w60, c1_n0_w61, c1_n0_w62, c1_n0_w63, c1_n0_w64, c1_n0_w65, c1_n0_w66, c1_n0_w67, c1_n0_w68, c1_n0_w69, c1_n0_w70, c1_n0_w71, c1_n0_w72, c1_n0_w73, c1_n0_w74, c1_n0_w75, c1_n0_w76, c1_n0_w77, c1_n0_w78, c1_n0_w79, c1_n0_w80, c1_n0_w81, c1_n0_w82, c1_n0_w83, c1_n0_w84, c1_n0_w85, c1_n0_w86, c1_n0_w87, c1_n0_w88, c1_n0_w89, c1_n0_w90, c1_n0_w91, c1_n0_w92, c1_n0_w93, c1_n0_w94, c1_n0_w95, c1_n0_w96, c1_n0_w97, c1_n0_w98, c1_n0_w99, c1_n0_w100, c1_n1_w1, c1_n1_w2, c1_n1_w3, c1_n1_w4, c1_n1_w5, c1_n1_w6, c1_n1_w7, c1_n1_w8, c1_n1_w9, c1_n1_w10, c1_n1_w11, c1_n1_w12, c1_n1_w13, c1_n1_w14, c1_n1_w15, c1_n1_w16, c1_n1_w17, c1_n1_w18, c1_n1_w19, c1_n1_w20, c1_n1_w21, c1_n1_w22, c1_n1_w23, c1_n1_w24, c1_n1_w25, c1_n1_w26, c1_n1_w27, c1_n1_w28, c1_n1_w29, c1_n1_w30, c1_n1_w31, c1_n1_w32, c1_n1_w33, c1_n1_w34, c1_n1_w35, c1_n1_w36, c1_n1_w37, c1_n1_w38, c1_n1_w39, c1_n1_w40, c1_n1_w41, c1_n1_w42, c1_n1_w43, c1_n1_w44, c1_n1_w45, c1_n1_w46, c1_n1_w47, c1_n1_w48, c1_n1_w49, c1_n1_w50, c1_n1_w51, c1_n1_w52, c1_n1_w53, c1_n1_w54, c1_n1_w55, c1_n1_w56, c1_n1_w57, c1_n1_w58, c1_n1_w59, c1_n1_w60, c1_n1_w61, c1_n1_w62, c1_n1_w63, c1_n1_w64, c1_n1_w65, c1_n1_w66, c1_n1_w67, c1_n1_w68, c1_n1_w69, c1_n1_w70, c1_n1_w71, c1_n1_w72, c1_n1_w73, c1_n1_w74, c1_n1_w75, c1_n1_w76, c1_n1_w77, c1_n1_w78, c1_n1_w79, c1_n1_w80, c1_n1_w81, c1_n1_w82, c1_n1_w83, c1_n1_w84, c1_n1_w85, c1_n1_w86, c1_n1_w87, c1_n1_w88, c1_n1_w89, c1_n1_w90, c1_n1_w91, c1_n1_w92, c1_n1_w93, c1_n1_w94, c1_n1_w95, c1_n1_w96, c1_n1_w97, c1_n1_w98, c1_n1_w99, c1_n1_w100, c1_n2_w1, c1_n2_w2, c1_n2_w3, c1_n2_w4, c1_n2_w5, c1_n2_w6, c1_n2_w7, c1_n2_w8, c1_n2_w9, c1_n2_w10, c1_n2_w11, c1_n2_w12, c1_n2_w13, c1_n2_w14, c1_n2_w15, c1_n2_w16, c1_n2_w17, c1_n2_w18, c1_n2_w19, c1_n2_w20, c1_n2_w21, c1_n2_w22, c1_n2_w23, c1_n2_w24, c1_n2_w25, c1_n2_w26, c1_n2_w27, c1_n2_w28, c1_n2_w29, c1_n2_w30, c1_n2_w31, c1_n2_w32, c1_n2_w33, c1_n2_w34, c1_n2_w35, c1_n2_w36, c1_n2_w37, c1_n2_w38, c1_n2_w39, c1_n2_w40, c1_n2_w41, c1_n2_w42, c1_n2_w43, c1_n2_w44, c1_n2_w45, c1_n2_w46, c1_n2_w47, c1_n2_w48, c1_n2_w49, c1_n2_w50, c1_n2_w51, c1_n2_w52, c1_n2_w53, c1_n2_w54, c1_n2_w55, c1_n2_w56, c1_n2_w57, c1_n2_w58, c1_n2_w59, c1_n2_w60, c1_n2_w61, c1_n2_w62, c1_n2_w63, c1_n2_w64, c1_n2_w65, c1_n2_w66, c1_n2_w67, c1_n2_w68, c1_n2_w69, c1_n2_w70, c1_n2_w71, c1_n2_w72, c1_n2_w73, c1_n2_w74, c1_n2_w75, c1_n2_w76, c1_n2_w77, c1_n2_w78, c1_n2_w79, c1_n2_w80, c1_n2_w81, c1_n2_w82, c1_n2_w83, c1_n2_w84, c1_n2_w85, c1_n2_w86, c1_n2_w87, c1_n2_w88, c1_n2_w89, c1_n2_w90, c1_n2_w91, c1_n2_w92, c1_n2_w93, c1_n2_w94, c1_n2_w95, c1_n2_w96, c1_n2_w97, c1_n2_w98, c1_n2_w99, c1_n2_w100, c1_n3_w1, c1_n3_w2, c1_n3_w3, c1_n3_w4, c1_n3_w5, c1_n3_w6, c1_n3_w7, c1_n3_w8, c1_n3_w9, c1_n3_w10, c1_n3_w11, c1_n3_w12, c1_n3_w13, c1_n3_w14, c1_n3_w15, c1_n3_w16, c1_n3_w17, c1_n3_w18, c1_n3_w19, c1_n3_w20, c1_n3_w21, c1_n3_w22, c1_n3_w23, c1_n3_w24, c1_n3_w25, c1_n3_w26, c1_n3_w27, c1_n3_w28, c1_n3_w29, c1_n3_w30, c1_n3_w31, c1_n3_w32, c1_n3_w33, c1_n3_w34, c1_n3_w35, c1_n3_w36, c1_n3_w37, c1_n3_w38, c1_n3_w39, c1_n3_w40, c1_n3_w41, c1_n3_w42, c1_n3_w43, c1_n3_w44, c1_n3_w45, c1_n3_w46, c1_n3_w47, c1_n3_w48, c1_n3_w49, c1_n3_w50, c1_n3_w51, c1_n3_w52, c1_n3_w53, c1_n3_w54, c1_n3_w55, c1_n3_w56, c1_n3_w57, c1_n3_w58, c1_n3_w59, c1_n3_w60, c1_n3_w61, c1_n3_w62, c1_n3_w63, c1_n3_w64, c1_n3_w65, c1_n3_w66, c1_n3_w67, c1_n3_w68, c1_n3_w69, c1_n3_w70, c1_n3_w71, c1_n3_w72, c1_n3_w73, c1_n3_w74, c1_n3_w75, c1_n3_w76, c1_n3_w77, c1_n3_w78, c1_n3_w79, c1_n3_w80, c1_n3_w81, c1_n3_w82, c1_n3_w83, c1_n3_w84, c1_n3_w85, c1_n3_w86, c1_n3_w87, c1_n3_w88, c1_n3_w89, c1_n3_w90, c1_n3_w91, c1_n3_w92, c1_n3_w93, c1_n3_w94, c1_n3_w95, c1_n3_w96, c1_n3_w97, c1_n3_w98, c1_n3_w99, c1_n3_w100, c1_n4_w1, c1_n4_w2, c1_n4_w3, c1_n4_w4, c1_n4_w5, c1_n4_w6, c1_n4_w7, c1_n4_w8, c1_n4_w9, c1_n4_w10, c1_n4_w11, c1_n4_w12, c1_n4_w13, c1_n4_w14, c1_n4_w15, c1_n4_w16, c1_n4_w17, c1_n4_w18, c1_n4_w19, c1_n4_w20, c1_n4_w21, c1_n4_w22, c1_n4_w23, c1_n4_w24, c1_n4_w25, c1_n4_w26, c1_n4_w27, c1_n4_w28, c1_n4_w29, c1_n4_w30, c1_n4_w31, c1_n4_w32, c1_n4_w33, c1_n4_w34, c1_n4_w35, c1_n4_w36, c1_n4_w37, c1_n4_w38, c1_n4_w39, c1_n4_w40, c1_n4_w41, c1_n4_w42, c1_n4_w43, c1_n4_w44, c1_n4_w45, c1_n4_w46, c1_n4_w47, c1_n4_w48, c1_n4_w49, c1_n4_w50, c1_n4_w51, c1_n4_w52, c1_n4_w53, c1_n4_w54, c1_n4_w55, c1_n4_w56, c1_n4_w57, c1_n4_w58, c1_n4_w59, c1_n4_w60, c1_n4_w61, c1_n4_w62, c1_n4_w63, c1_n4_w64, c1_n4_w65, c1_n4_w66, c1_n4_w67, c1_n4_w68, c1_n4_w69, c1_n4_w70, c1_n4_w71, c1_n4_w72, c1_n4_w73, c1_n4_w74, c1_n4_w75, c1_n4_w76, c1_n4_w77, c1_n4_w78, c1_n4_w79, c1_n4_w80, c1_n4_w81, c1_n4_w82, c1_n4_w83, c1_n4_w84, c1_n4_w85, c1_n4_w86, c1_n4_w87, c1_n4_w88, c1_n4_w89, c1_n4_w90, c1_n4_w91, c1_n4_w92, c1_n4_w93, c1_n4_w94, c1_n4_w95, c1_n4_w96, c1_n4_w97, c1_n4_w98, c1_n4_w99, c1_n4_w100, c1_n5_w1, c1_n5_w2, c1_n5_w3, c1_n5_w4, c1_n5_w5, c1_n5_w6, c1_n5_w7, c1_n5_w8, c1_n5_w9, c1_n5_w10, c1_n5_w11, c1_n5_w12, c1_n5_w13, c1_n5_w14, c1_n5_w15, c1_n5_w16, c1_n5_w17, c1_n5_w18, c1_n5_w19, c1_n5_w20, c1_n5_w21, c1_n5_w22, c1_n5_w23, c1_n5_w24, c1_n5_w25, c1_n5_w26, c1_n5_w27, c1_n5_w28, c1_n5_w29, c1_n5_w30, c1_n5_w31, c1_n5_w32, c1_n5_w33, c1_n5_w34, c1_n5_w35, c1_n5_w36, c1_n5_w37, c1_n5_w38, c1_n5_w39, c1_n5_w40, c1_n5_w41, c1_n5_w42, c1_n5_w43, c1_n5_w44, c1_n5_w45, c1_n5_w46, c1_n5_w47, c1_n5_w48, c1_n5_w49, c1_n5_w50, c1_n5_w51, c1_n5_w52, c1_n5_w53, c1_n5_w54, c1_n5_w55, c1_n5_w56, c1_n5_w57, c1_n5_w58, c1_n5_w59, c1_n5_w60, c1_n5_w61, c1_n5_w62, c1_n5_w63, c1_n5_w64, c1_n5_w65, c1_n5_w66, c1_n5_w67, c1_n5_w68, c1_n5_w69, c1_n5_w70, c1_n5_w71, c1_n5_w72, c1_n5_w73, c1_n5_w74, c1_n5_w75, c1_n5_w76, c1_n5_w77, c1_n5_w78, c1_n5_w79, c1_n5_w80, c1_n5_w81, c1_n5_w82, c1_n5_w83, c1_n5_w84, c1_n5_w85, c1_n5_w86, c1_n5_w87, c1_n5_w88, c1_n5_w89, c1_n5_w90, c1_n5_w91, c1_n5_w92, c1_n5_w93, c1_n5_w94, c1_n5_w95, c1_n5_w96, c1_n5_w97, c1_n5_w98, c1_n5_w99, c1_n5_w100, c1_n6_w1, c1_n6_w2, c1_n6_w3, c1_n6_w4, c1_n6_w5, c1_n6_w6, c1_n6_w7, c1_n6_w8, c1_n6_w9, c1_n6_w10, c1_n6_w11, c1_n6_w12, c1_n6_w13, c1_n6_w14, c1_n6_w15, c1_n6_w16, c1_n6_w17, c1_n6_w18, c1_n6_w19, c1_n6_w20, c1_n6_w21, c1_n6_w22, c1_n6_w23, c1_n6_w24, c1_n6_w25, c1_n6_w26, c1_n6_w27, c1_n6_w28, c1_n6_w29, c1_n6_w30, c1_n6_w31, c1_n6_w32, c1_n6_w33, c1_n6_w34, c1_n6_w35, c1_n6_w36, c1_n6_w37, c1_n6_w38, c1_n6_w39, c1_n6_w40, c1_n6_w41, c1_n6_w42, c1_n6_w43, c1_n6_w44, c1_n6_w45, c1_n6_w46, c1_n6_w47, c1_n6_w48, c1_n6_w49, c1_n6_w50, c1_n6_w51, c1_n6_w52, c1_n6_w53, c1_n6_w54, c1_n6_w55, c1_n6_w56, c1_n6_w57, c1_n6_w58, c1_n6_w59, c1_n6_w60, c1_n6_w61, c1_n6_w62, c1_n6_w63, c1_n6_w64, c1_n6_w65, c1_n6_w66, c1_n6_w67, c1_n6_w68, c1_n6_w69, c1_n6_w70, c1_n6_w71, c1_n6_w72, c1_n6_w73, c1_n6_w74, c1_n6_w75, c1_n6_w76, c1_n6_w77, c1_n6_w78, c1_n6_w79, c1_n6_w80, c1_n6_w81, c1_n6_w82, c1_n6_w83, c1_n6_w84, c1_n6_w85, c1_n6_w86, c1_n6_w87, c1_n6_w88, c1_n6_w89, c1_n6_w90, c1_n6_w91, c1_n6_w92, c1_n6_w93, c1_n6_w94, c1_n6_w95, c1_n6_w96, c1_n6_w97, c1_n6_w98, c1_n6_w99, c1_n6_w100, c1_n7_w1, c1_n7_w2, c1_n7_w3, c1_n7_w4, c1_n7_w5, c1_n7_w6, c1_n7_w7, c1_n7_w8, c1_n7_w9, c1_n7_w10, c1_n7_w11, c1_n7_w12, c1_n7_w13, c1_n7_w14, c1_n7_w15, c1_n7_w16, c1_n7_w17, c1_n7_w18, c1_n7_w19, c1_n7_w20, c1_n7_w21, c1_n7_w22, c1_n7_w23, c1_n7_w24, c1_n7_w25, c1_n7_w26, c1_n7_w27, c1_n7_w28, c1_n7_w29, c1_n7_w30, c1_n7_w31, c1_n7_w32, c1_n7_w33, c1_n7_w34, c1_n7_w35, c1_n7_w36, c1_n7_w37, c1_n7_w38, c1_n7_w39, c1_n7_w40, c1_n7_w41, c1_n7_w42, c1_n7_w43, c1_n7_w44, c1_n7_w45, c1_n7_w46, c1_n7_w47, c1_n7_w48, c1_n7_w49, c1_n7_w50, c1_n7_w51, c1_n7_w52, c1_n7_w53, c1_n7_w54, c1_n7_w55, c1_n7_w56, c1_n7_w57, c1_n7_w58, c1_n7_w59, c1_n7_w60, c1_n7_w61, c1_n7_w62, c1_n7_w63, c1_n7_w64, c1_n7_w65, c1_n7_w66, c1_n7_w67, c1_n7_w68, c1_n7_w69, c1_n7_w70, c1_n7_w71, c1_n7_w72, c1_n7_w73, c1_n7_w74, c1_n7_w75, c1_n7_w76, c1_n7_w77, c1_n7_w78, c1_n7_w79, c1_n7_w80, c1_n7_w81, c1_n7_w82, c1_n7_w83, c1_n7_w84, c1_n7_w85, c1_n7_w86, c1_n7_w87, c1_n7_w88, c1_n7_w89, c1_n7_w90, c1_n7_w91, c1_n7_w92, c1_n7_w93, c1_n7_w94, c1_n7_w95, c1_n7_w96, c1_n7_w97, c1_n7_w98, c1_n7_w99, c1_n7_w100, c1_n8_w1, c1_n8_w2, c1_n8_w3, c1_n8_w4, c1_n8_w5, c1_n8_w6, c1_n8_w7, c1_n8_w8, c1_n8_w9, c1_n8_w10, c1_n8_w11, c1_n8_w12, c1_n8_w13, c1_n8_w14, c1_n8_w15, c1_n8_w16, c1_n8_w17, c1_n8_w18, c1_n8_w19, c1_n8_w20, c1_n8_w21, c1_n8_w22, c1_n8_w23, c1_n8_w24, c1_n8_w25, c1_n8_w26, c1_n8_w27, c1_n8_w28, c1_n8_w29, c1_n8_w30, c1_n8_w31, c1_n8_w32, c1_n8_w33, c1_n8_w34, c1_n8_w35, c1_n8_w36, c1_n8_w37, c1_n8_w38, c1_n8_w39, c1_n8_w40, c1_n8_w41, c1_n8_w42, c1_n8_w43, c1_n8_w44, c1_n8_w45, c1_n8_w46, c1_n8_w47, c1_n8_w48, c1_n8_w49, c1_n8_w50, c1_n8_w51, c1_n8_w52, c1_n8_w53, c1_n8_w54, c1_n8_w55, c1_n8_w56, c1_n8_w57, c1_n8_w58, c1_n8_w59, c1_n8_w60, c1_n8_w61, c1_n8_w62, c1_n8_w63, c1_n8_w64, c1_n8_w65, c1_n8_w66, c1_n8_w67, c1_n8_w68, c1_n8_w69, c1_n8_w70, c1_n8_w71, c1_n8_w72, c1_n8_w73, c1_n8_w74, c1_n8_w75, c1_n8_w76, c1_n8_w77, c1_n8_w78, c1_n8_w79, c1_n8_w80, c1_n8_w81, c1_n8_w82, c1_n8_w83, c1_n8_w84, c1_n8_w85, c1_n8_w86, c1_n8_w87, c1_n8_w88, c1_n8_w89, c1_n8_w90, c1_n8_w91, c1_n8_w92, c1_n8_w93, c1_n8_w94, c1_n8_w95, c1_n8_w96, c1_n8_w97, c1_n8_w98, c1_n8_w99, c1_n8_w100, c1_n9_w1, c1_n9_w2, c1_n9_w3, c1_n9_w4, c1_n9_w5, c1_n9_w6, c1_n9_w7, c1_n9_w8, c1_n9_w9, c1_n9_w10, c1_n9_w11, c1_n9_w12, c1_n9_w13, c1_n9_w14, c1_n9_w15, c1_n9_w16, c1_n9_w17, c1_n9_w18, c1_n9_w19, c1_n9_w20, c1_n9_w21, c1_n9_w22, c1_n9_w23, c1_n9_w24, c1_n9_w25, c1_n9_w26, c1_n9_w27, c1_n9_w28, c1_n9_w29, c1_n9_w30, c1_n9_w31, c1_n9_w32, c1_n9_w33, c1_n9_w34, c1_n9_w35, c1_n9_w36, c1_n9_w37, c1_n9_w38, c1_n9_w39, c1_n9_w40, c1_n9_w41, c1_n9_w42, c1_n9_w43, c1_n9_w44, c1_n9_w45, c1_n9_w46, c1_n9_w47, c1_n9_w48, c1_n9_w49, c1_n9_w50, c1_n9_w51, c1_n9_w52, c1_n9_w53, c1_n9_w54, c1_n9_w55, c1_n9_w56, c1_n9_w57, c1_n9_w58, c1_n9_w59, c1_n9_w60, c1_n9_w61, c1_n9_w62, c1_n9_w63, c1_n9_w64, c1_n9_w65, c1_n9_w66, c1_n9_w67, c1_n9_w68, c1_n9_w69, c1_n9_w70, c1_n9_w71, c1_n9_w72, c1_n9_w73, c1_n9_w74, c1_n9_w75, c1_n9_w76, c1_n9_w77, c1_n9_w78, c1_n9_w79, c1_n9_w80, c1_n9_w81, c1_n9_w82, c1_n9_w83, c1_n9_w84, c1_n9_w85, c1_n9_w86, c1_n9_w87, c1_n9_w88, c1_n9_w89, c1_n9_w90, c1_n9_w91, c1_n9_w92, c1_n9_w93, c1_n9_w94, c1_n9_w95, c1_n9_w96, c1_n9_w97, c1_n9_w98, c1_n9_w99, c1_n9_w100, c1_n10_w1, c1_n10_w2, c1_n10_w3, c1_n10_w4, c1_n10_w5, c1_n10_w6, c1_n10_w7, c1_n10_w8, c1_n10_w9, c1_n10_w10, c1_n10_w11, c1_n10_w12, c1_n10_w13, c1_n10_w14, c1_n10_w15, c1_n10_w16, c1_n10_w17, c1_n10_w18, c1_n10_w19, c1_n10_w20, c1_n10_w21, c1_n10_w22, c1_n10_w23, c1_n10_w24, c1_n10_w25, c1_n10_w26, c1_n10_w27, c1_n10_w28, c1_n10_w29, c1_n10_w30, c1_n10_w31, c1_n10_w32, c1_n10_w33, c1_n10_w34, c1_n10_w35, c1_n10_w36, c1_n10_w37, c1_n10_w38, c1_n10_w39, c1_n10_w40, c1_n10_w41, c1_n10_w42, c1_n10_w43, c1_n10_w44, c1_n10_w45, c1_n10_w46, c1_n10_w47, c1_n10_w48, c1_n10_w49, c1_n10_w50, c1_n10_w51, c1_n10_w52, c1_n10_w53, c1_n10_w54, c1_n10_w55, c1_n10_w56, c1_n10_w57, c1_n10_w58, c1_n10_w59, c1_n10_w60, c1_n10_w61, c1_n10_w62, c1_n10_w63, c1_n10_w64, c1_n10_w65, c1_n10_w66, c1_n10_w67, c1_n10_w68, c1_n10_w69, c1_n10_w70, c1_n10_w71, c1_n10_w72, c1_n10_w73, c1_n10_w74, c1_n10_w75, c1_n10_w76, c1_n10_w77, c1_n10_w78, c1_n10_w79, c1_n10_w80, c1_n10_w81, c1_n10_w82, c1_n10_w83, c1_n10_w84, c1_n10_w85, c1_n10_w86, c1_n10_w87, c1_n10_w88, c1_n10_w89, c1_n10_w90, c1_n10_w91, c1_n10_w92, c1_n10_w93, c1_n10_w94, c1_n10_w95, c1_n10_w96, c1_n10_w97, c1_n10_w98, c1_n10_w99, c1_n10_w100, c1_n11_w1, c1_n11_w2, c1_n11_w3, c1_n11_w4, c1_n11_w5, c1_n11_w6, c1_n11_w7, c1_n11_w8, c1_n11_w9, c1_n11_w10, c1_n11_w11, c1_n11_w12, c1_n11_w13, c1_n11_w14, c1_n11_w15, c1_n11_w16, c1_n11_w17, c1_n11_w18, c1_n11_w19, c1_n11_w20, c1_n11_w21, c1_n11_w22, c1_n11_w23, c1_n11_w24, c1_n11_w25, c1_n11_w26, c1_n11_w27, c1_n11_w28, c1_n11_w29, c1_n11_w30, c1_n11_w31, c1_n11_w32, c1_n11_w33, c1_n11_w34, c1_n11_w35, c1_n11_w36, c1_n11_w37, c1_n11_w38, c1_n11_w39, c1_n11_w40, c1_n11_w41, c1_n11_w42, c1_n11_w43, c1_n11_w44, c1_n11_w45, c1_n11_w46, c1_n11_w47, c1_n11_w48, c1_n11_w49, c1_n11_w50, c1_n11_w51, c1_n11_w52, c1_n11_w53, c1_n11_w54, c1_n11_w55, c1_n11_w56, c1_n11_w57, c1_n11_w58, c1_n11_w59, c1_n11_w60, c1_n11_w61, c1_n11_w62, c1_n11_w63, c1_n11_w64, c1_n11_w65, c1_n11_w66, c1_n11_w67, c1_n11_w68, c1_n11_w69, c1_n11_w70, c1_n11_w71, c1_n11_w72, c1_n11_w73, c1_n11_w74, c1_n11_w75, c1_n11_w76, c1_n11_w77, c1_n11_w78, c1_n11_w79, c1_n11_w80, c1_n11_w81, c1_n11_w82, c1_n11_w83, c1_n11_w84, c1_n11_w85, c1_n11_w86, c1_n11_w87, c1_n11_w88, c1_n11_w89, c1_n11_w90, c1_n11_w91, c1_n11_w92, c1_n11_w93, c1_n11_w94, c1_n11_w95, c1_n11_w96, c1_n11_w97, c1_n11_w98, c1_n11_w99, c1_n11_w100, c1_n12_w1, c1_n12_w2, c1_n12_w3, c1_n12_w4, c1_n12_w5, c1_n12_w6, c1_n12_w7, c1_n12_w8, c1_n12_w9, c1_n12_w10, c1_n12_w11, c1_n12_w12, c1_n12_w13, c1_n12_w14, c1_n12_w15, c1_n12_w16, c1_n12_w17, c1_n12_w18, c1_n12_w19, c1_n12_w20, c1_n12_w21, c1_n12_w22, c1_n12_w23, c1_n12_w24, c1_n12_w25, c1_n12_w26, c1_n12_w27, c1_n12_w28, c1_n12_w29, c1_n12_w30, c1_n12_w31, c1_n12_w32, c1_n12_w33, c1_n12_w34, c1_n12_w35, c1_n12_w36, c1_n12_w37, c1_n12_w38, c1_n12_w39, c1_n12_w40, c1_n12_w41, c1_n12_w42, c1_n12_w43, c1_n12_w44, c1_n12_w45, c1_n12_w46, c1_n12_w47, c1_n12_w48, c1_n12_w49, c1_n12_w50, c1_n12_w51, c1_n12_w52, c1_n12_w53, c1_n12_w54, c1_n12_w55, c1_n12_w56, c1_n12_w57, c1_n12_w58, c1_n12_w59, c1_n12_w60, c1_n12_w61, c1_n12_w62, c1_n12_w63, c1_n12_w64, c1_n12_w65, c1_n12_w66, c1_n12_w67, c1_n12_w68, c1_n12_w69, c1_n12_w70, c1_n12_w71, c1_n12_w72, c1_n12_w73, c1_n12_w74, c1_n12_w75, c1_n12_w76, c1_n12_w77, c1_n12_w78, c1_n12_w79, c1_n12_w80, c1_n12_w81, c1_n12_w82, c1_n12_w83, c1_n12_w84, c1_n12_w85, c1_n12_w86, c1_n12_w87, c1_n12_w88, c1_n12_w89, c1_n12_w90, c1_n12_w91, c1_n12_w92, c1_n12_w93, c1_n12_w94, c1_n12_w95, c1_n12_w96, c1_n12_w97, c1_n12_w98, c1_n12_w99, c1_n12_w100, c1_n13_w1, c1_n13_w2, c1_n13_w3, c1_n13_w4, c1_n13_w5, c1_n13_w6, c1_n13_w7, c1_n13_w8, c1_n13_w9, c1_n13_w10, c1_n13_w11, c1_n13_w12, c1_n13_w13, c1_n13_w14, c1_n13_w15, c1_n13_w16, c1_n13_w17, c1_n13_w18, c1_n13_w19, c1_n13_w20, c1_n13_w21, c1_n13_w22, c1_n13_w23, c1_n13_w24, c1_n13_w25, c1_n13_w26, c1_n13_w27, c1_n13_w28, c1_n13_w29, c1_n13_w30, c1_n13_w31, c1_n13_w32, c1_n13_w33, c1_n13_w34, c1_n13_w35, c1_n13_w36, c1_n13_w37, c1_n13_w38, c1_n13_w39, c1_n13_w40, c1_n13_w41, c1_n13_w42, c1_n13_w43, c1_n13_w44, c1_n13_w45, c1_n13_w46, c1_n13_w47, c1_n13_w48, c1_n13_w49, c1_n13_w50, c1_n13_w51, c1_n13_w52, c1_n13_w53, c1_n13_w54, c1_n13_w55, c1_n13_w56, c1_n13_w57, c1_n13_w58, c1_n13_w59, c1_n13_w60, c1_n13_w61, c1_n13_w62, c1_n13_w63, c1_n13_w64, c1_n13_w65, c1_n13_w66, c1_n13_w67, c1_n13_w68, c1_n13_w69, c1_n13_w70, c1_n13_w71, c1_n13_w72, c1_n13_w73, c1_n13_w74, c1_n13_w75, c1_n13_w76, c1_n13_w77, c1_n13_w78, c1_n13_w79, c1_n13_w80, c1_n13_w81, c1_n13_w82, c1_n13_w83, c1_n13_w84, c1_n13_w85, c1_n13_w86, c1_n13_w87, c1_n13_w88, c1_n13_w89, c1_n13_w90, c1_n13_w91, c1_n13_w92, c1_n13_w93, c1_n13_w94, c1_n13_w95, c1_n13_w96, c1_n13_w97, c1_n13_w98, c1_n13_w99, c1_n13_w100, c1_n14_w1, c1_n14_w2, c1_n14_w3, c1_n14_w4, c1_n14_w5, c1_n14_w6, c1_n14_w7, c1_n14_w8, c1_n14_w9, c1_n14_w10, c1_n14_w11, c1_n14_w12, c1_n14_w13, c1_n14_w14, c1_n14_w15, c1_n14_w16, c1_n14_w17, c1_n14_w18, c1_n14_w19, c1_n14_w20, c1_n14_w21, c1_n14_w22, c1_n14_w23, c1_n14_w24, c1_n14_w25, c1_n14_w26, c1_n14_w27, c1_n14_w28, c1_n14_w29, c1_n14_w30, c1_n14_w31, c1_n14_w32, c1_n14_w33, c1_n14_w34, c1_n14_w35, c1_n14_w36, c1_n14_w37, c1_n14_w38, c1_n14_w39, c1_n14_w40, c1_n14_w41, c1_n14_w42, c1_n14_w43, c1_n14_w44, c1_n14_w45, c1_n14_w46, c1_n14_w47, c1_n14_w48, c1_n14_w49, c1_n14_w50, c1_n14_w51, c1_n14_w52, c1_n14_w53, c1_n14_w54, c1_n14_w55, c1_n14_w56, c1_n14_w57, c1_n14_w58, c1_n14_w59, c1_n14_w60, c1_n14_w61, c1_n14_w62, c1_n14_w63, c1_n14_w64, c1_n14_w65, c1_n14_w66, c1_n14_w67, c1_n14_w68, c1_n14_w69, c1_n14_w70, c1_n14_w71, c1_n14_w72, c1_n14_w73, c1_n14_w74, c1_n14_w75, c1_n14_w76, c1_n14_w77, c1_n14_w78, c1_n14_w79, c1_n14_w80, c1_n14_w81, c1_n14_w82, c1_n14_w83, c1_n14_w84, c1_n14_w85, c1_n14_w86, c1_n14_w87, c1_n14_w88, c1_n14_w89, c1_n14_w90, c1_n14_w91, c1_n14_w92, c1_n14_w93, c1_n14_w94, c1_n14_w95, c1_n14_w96, c1_n14_w97, c1_n14_w98, c1_n14_w99, c1_n14_w100, c1_n15_w1, c1_n15_w2, c1_n15_w3, c1_n15_w4, c1_n15_w5, c1_n15_w6, c1_n15_w7, c1_n15_w8, c1_n15_w9, c1_n15_w10, c1_n15_w11, c1_n15_w12, c1_n15_w13, c1_n15_w14, c1_n15_w15, c1_n15_w16, c1_n15_w17, c1_n15_w18, c1_n15_w19, c1_n15_w20, c1_n15_w21, c1_n15_w22, c1_n15_w23, c1_n15_w24, c1_n15_w25, c1_n15_w26, c1_n15_w27, c1_n15_w28, c1_n15_w29, c1_n15_w30, c1_n15_w31, c1_n15_w32, c1_n15_w33, c1_n15_w34, c1_n15_w35, c1_n15_w36, c1_n15_w37, c1_n15_w38, c1_n15_w39, c1_n15_w40, c1_n15_w41, c1_n15_w42, c1_n15_w43, c1_n15_w44, c1_n15_w45, c1_n15_w46, c1_n15_w47, c1_n15_w48, c1_n15_w49, c1_n15_w50, c1_n15_w51, c1_n15_w52, c1_n15_w53, c1_n15_w54, c1_n15_w55, c1_n15_w56, c1_n15_w57, c1_n15_w58, c1_n15_w59, c1_n15_w60, c1_n15_w61, c1_n15_w62, c1_n15_w63, c1_n15_w64, c1_n15_w65, c1_n15_w66, c1_n15_w67, c1_n15_w68, c1_n15_w69, c1_n15_w70, c1_n15_w71, c1_n15_w72, c1_n15_w73, c1_n15_w74, c1_n15_w75, c1_n15_w76, c1_n15_w77, c1_n15_w78, c1_n15_w79, c1_n15_w80, c1_n15_w81, c1_n15_w82, c1_n15_w83, c1_n15_w84, c1_n15_w85, c1_n15_w86, c1_n15_w87, c1_n15_w88, c1_n15_w89, c1_n15_w90, c1_n15_w91, c1_n15_w92, c1_n15_w93, c1_n15_w94, c1_n15_w95, c1_n15_w96, c1_n15_w97, c1_n15_w98, c1_n15_w99, c1_n15_w100, c1_n16_w1, c1_n16_w2, c1_n16_w3, c1_n16_w4, c1_n16_w5, c1_n16_w6, c1_n16_w7, c1_n16_w8, c1_n16_w9, c1_n16_w10, c1_n16_w11, c1_n16_w12, c1_n16_w13, c1_n16_w14, c1_n16_w15, c1_n16_w16, c1_n16_w17, c1_n16_w18, c1_n16_w19, c1_n16_w20, c1_n16_w21, c1_n16_w22, c1_n16_w23, c1_n16_w24, c1_n16_w25, c1_n16_w26, c1_n16_w27, c1_n16_w28, c1_n16_w29, c1_n16_w30, c1_n16_w31, c1_n16_w32, c1_n16_w33, c1_n16_w34, c1_n16_w35, c1_n16_w36, c1_n16_w37, c1_n16_w38, c1_n16_w39, c1_n16_w40, c1_n16_w41, c1_n16_w42, c1_n16_w43, c1_n16_w44, c1_n16_w45, c1_n16_w46, c1_n16_w47, c1_n16_w48, c1_n16_w49, c1_n16_w50, c1_n16_w51, c1_n16_w52, c1_n16_w53, c1_n16_w54, c1_n16_w55, c1_n16_w56, c1_n16_w57, c1_n16_w58, c1_n16_w59, c1_n16_w60, c1_n16_w61, c1_n16_w62, c1_n16_w63, c1_n16_w64, c1_n16_w65, c1_n16_w66, c1_n16_w67, c1_n16_w68, c1_n16_w69, c1_n16_w70, c1_n16_w71, c1_n16_w72, c1_n16_w73, c1_n16_w74, c1_n16_w75, c1_n16_w76, c1_n16_w77, c1_n16_w78, c1_n16_w79, c1_n16_w80, c1_n16_w81, c1_n16_w82, c1_n16_w83, c1_n16_w84, c1_n16_w85, c1_n16_w86, c1_n16_w87, c1_n16_w88, c1_n16_w89, c1_n16_w90, c1_n16_w91, c1_n16_w92, c1_n16_w93, c1_n16_w94, c1_n16_w95, c1_n16_w96, c1_n16_w97, c1_n16_w98, c1_n16_w99, c1_n16_w100, c1_n17_w1, c1_n17_w2, c1_n17_w3, c1_n17_w4, c1_n17_w5, c1_n17_w6, c1_n17_w7, c1_n17_w8, c1_n17_w9, c1_n17_w10, c1_n17_w11, c1_n17_w12, c1_n17_w13, c1_n17_w14, c1_n17_w15, c1_n17_w16, c1_n17_w17, c1_n17_w18, c1_n17_w19, c1_n17_w20, c1_n17_w21, c1_n17_w22, c1_n17_w23, c1_n17_w24, c1_n17_w25, c1_n17_w26, c1_n17_w27, c1_n17_w28, c1_n17_w29, c1_n17_w30, c1_n17_w31, c1_n17_w32, c1_n17_w33, c1_n17_w34, c1_n17_w35, c1_n17_w36, c1_n17_w37, c1_n17_w38, c1_n17_w39, c1_n17_w40, c1_n17_w41, c1_n17_w42, c1_n17_w43, c1_n17_w44, c1_n17_w45, c1_n17_w46, c1_n17_w47, c1_n17_w48, c1_n17_w49, c1_n17_w50, c1_n17_w51, c1_n17_w52, c1_n17_w53, c1_n17_w54, c1_n17_w55, c1_n17_w56, c1_n17_w57, c1_n17_w58, c1_n17_w59, c1_n17_w60, c1_n17_w61, c1_n17_w62, c1_n17_w63, c1_n17_w64, c1_n17_w65, c1_n17_w66, c1_n17_w67, c1_n17_w68, c1_n17_w69, c1_n17_w70, c1_n17_w71, c1_n17_w72, c1_n17_w73, c1_n17_w74, c1_n17_w75, c1_n17_w76, c1_n17_w77, c1_n17_w78, c1_n17_w79, c1_n17_w80, c1_n17_w81, c1_n17_w82, c1_n17_w83, c1_n17_w84, c1_n17_w85, c1_n17_w86, c1_n17_w87, c1_n17_w88, c1_n17_w89, c1_n17_w90, c1_n17_w91, c1_n17_w92, c1_n17_w93, c1_n17_w94, c1_n17_w95, c1_n17_w96, c1_n17_w97, c1_n17_w98, c1_n17_w99, c1_n17_w100, c1_n18_w1, c1_n18_w2, c1_n18_w3, c1_n18_w4, c1_n18_w5, c1_n18_w6, c1_n18_w7, c1_n18_w8, c1_n18_w9, c1_n18_w10, c1_n18_w11, c1_n18_w12, c1_n18_w13, c1_n18_w14, c1_n18_w15, c1_n18_w16, c1_n18_w17, c1_n18_w18, c1_n18_w19, c1_n18_w20, c1_n18_w21, c1_n18_w22, c1_n18_w23, c1_n18_w24, c1_n18_w25, c1_n18_w26, c1_n18_w27, c1_n18_w28, c1_n18_w29, c1_n18_w30, c1_n18_w31, c1_n18_w32, c1_n18_w33, c1_n18_w34, c1_n18_w35, c1_n18_w36, c1_n18_w37, c1_n18_w38, c1_n18_w39, c1_n18_w40, c1_n18_w41, c1_n18_w42, c1_n18_w43, c1_n18_w44, c1_n18_w45, c1_n18_w46, c1_n18_w47, c1_n18_w48, c1_n18_w49, c1_n18_w50, c1_n18_w51, c1_n18_w52, c1_n18_w53, c1_n18_w54, c1_n18_w55, c1_n18_w56, c1_n18_w57, c1_n18_w58, c1_n18_w59, c1_n18_w60, c1_n18_w61, c1_n18_w62, c1_n18_w63, c1_n18_w64, c1_n18_w65, c1_n18_w66, c1_n18_w67, c1_n18_w68, c1_n18_w69, c1_n18_w70, c1_n18_w71, c1_n18_w72, c1_n18_w73, c1_n18_w74, c1_n18_w75, c1_n18_w76, c1_n18_w77, c1_n18_w78, c1_n18_w79, c1_n18_w80, c1_n18_w81, c1_n18_w82, c1_n18_w83, c1_n18_w84, c1_n18_w85, c1_n18_w86, c1_n18_w87, c1_n18_w88, c1_n18_w89, c1_n18_w90, c1_n18_w91, c1_n18_w92, c1_n18_w93, c1_n18_w94, c1_n18_w95, c1_n18_w96, c1_n18_w97, c1_n18_w98, c1_n18_w99, c1_n18_w100, c1_n19_w1, c1_n19_w2, c1_n19_w3, c1_n19_w4, c1_n19_w5, c1_n19_w6, c1_n19_w7, c1_n19_w8, c1_n19_w9, c1_n19_w10, c1_n19_w11, c1_n19_w12, c1_n19_w13, c1_n19_w14, c1_n19_w15, c1_n19_w16, c1_n19_w17, c1_n19_w18, c1_n19_w19, c1_n19_w20, c1_n19_w21, c1_n19_w22, c1_n19_w23, c1_n19_w24, c1_n19_w25, c1_n19_w26, c1_n19_w27, c1_n19_w28, c1_n19_w29, c1_n19_w30, c1_n19_w31, c1_n19_w32, c1_n19_w33, c1_n19_w34, c1_n19_w35, c1_n19_w36, c1_n19_w37, c1_n19_w38, c1_n19_w39, c1_n19_w40, c1_n19_w41, c1_n19_w42, c1_n19_w43, c1_n19_w44, c1_n19_w45, c1_n19_w46, c1_n19_w47, c1_n19_w48, c1_n19_w49, c1_n19_w50, c1_n19_w51, c1_n19_w52, c1_n19_w53, c1_n19_w54, c1_n19_w55, c1_n19_w56, c1_n19_w57, c1_n19_w58, c1_n19_w59, c1_n19_w60, c1_n19_w61, c1_n19_w62, c1_n19_w63, c1_n19_w64, c1_n19_w65, c1_n19_w66, c1_n19_w67, c1_n19_w68, c1_n19_w69, c1_n19_w70, c1_n19_w71, c1_n19_w72, c1_n19_w73, c1_n19_w74, c1_n19_w75, c1_n19_w76, c1_n19_w77, c1_n19_w78, c1_n19_w79, c1_n19_w80, c1_n19_w81, c1_n19_w82, c1_n19_w83, c1_n19_w84, c1_n19_w85, c1_n19_w86, c1_n19_w87, c1_n19_w88, c1_n19_w89, c1_n19_w90, c1_n19_w91, c1_n19_w92, c1_n19_w93, c1_n19_w94, c1_n19_w95, c1_n19_w96, c1_n19_w97, c1_n19_w98, c1_n19_w99, c1_n19_w100, c1_n20_w1, c1_n20_w2, c1_n20_w3, c1_n20_w4, c1_n20_w5, c1_n20_w6, c1_n20_w7, c1_n20_w8, c1_n20_w9, c1_n20_w10, c1_n20_w11, c1_n20_w12, c1_n20_w13, c1_n20_w14, c1_n20_w15, c1_n20_w16, c1_n20_w17, c1_n20_w18, c1_n20_w19, c1_n20_w20, c1_n20_w21, c1_n20_w22, c1_n20_w23, c1_n20_w24, c1_n20_w25, c1_n20_w26, c1_n20_w27, c1_n20_w28, c1_n20_w29, c1_n20_w30, c1_n20_w31, c1_n20_w32, c1_n20_w33, c1_n20_w34, c1_n20_w35, c1_n20_w36, c1_n20_w37, c1_n20_w38, c1_n20_w39, c1_n20_w40, c1_n20_w41, c1_n20_w42, c1_n20_w43, c1_n20_w44, c1_n20_w45, c1_n20_w46, c1_n20_w47, c1_n20_w48, c1_n20_w49, c1_n20_w50, c1_n20_w51, c1_n20_w52, c1_n20_w53, c1_n20_w54, c1_n20_w55, c1_n20_w56, c1_n20_w57, c1_n20_w58, c1_n20_w59, c1_n20_w60, c1_n20_w61, c1_n20_w62, c1_n20_w63, c1_n20_w64, c1_n20_w65, c1_n20_w66, c1_n20_w67, c1_n20_w68, c1_n20_w69, c1_n20_w70, c1_n20_w71, c1_n20_w72, c1_n20_w73, c1_n20_w74, c1_n20_w75, c1_n20_w76, c1_n20_w77, c1_n20_w78, c1_n20_w79, c1_n20_w80, c1_n20_w81, c1_n20_w82, c1_n20_w83, c1_n20_w84, c1_n20_w85, c1_n20_w86, c1_n20_w87, c1_n20_w88, c1_n20_w89, c1_n20_w90, c1_n20_w91, c1_n20_w92, c1_n20_w93, c1_n20_w94, c1_n20_w95, c1_n20_w96, c1_n20_w97, c1_n20_w98, c1_n20_w99, c1_n20_w100, c1_n21_w1, c1_n21_w2, c1_n21_w3, c1_n21_w4, c1_n21_w5, c1_n21_w6, c1_n21_w7, c1_n21_w8, c1_n21_w9, c1_n21_w10, c1_n21_w11, c1_n21_w12, c1_n21_w13, c1_n21_w14, c1_n21_w15, c1_n21_w16, c1_n21_w17, c1_n21_w18, c1_n21_w19, c1_n21_w20, c1_n21_w21, c1_n21_w22, c1_n21_w23, c1_n21_w24, c1_n21_w25, c1_n21_w26, c1_n21_w27, c1_n21_w28, c1_n21_w29, c1_n21_w30, c1_n21_w31, c1_n21_w32, c1_n21_w33, c1_n21_w34, c1_n21_w35, c1_n21_w36, c1_n21_w37, c1_n21_w38, c1_n21_w39, c1_n21_w40, c1_n21_w41, c1_n21_w42, c1_n21_w43, c1_n21_w44, c1_n21_w45, c1_n21_w46, c1_n21_w47, c1_n21_w48, c1_n21_w49, c1_n21_w50, c1_n21_w51, c1_n21_w52, c1_n21_w53, c1_n21_w54, c1_n21_w55, c1_n21_w56, c1_n21_w57, c1_n21_w58, c1_n21_w59, c1_n21_w60, c1_n21_w61, c1_n21_w62, c1_n21_w63, c1_n21_w64, c1_n21_w65, c1_n21_w66, c1_n21_w67, c1_n21_w68, c1_n21_w69, c1_n21_w70, c1_n21_w71, c1_n21_w72, c1_n21_w73, c1_n21_w74, c1_n21_w75, c1_n21_w76, c1_n21_w77, c1_n21_w78, c1_n21_w79, c1_n21_w80, c1_n21_w81, c1_n21_w82, c1_n21_w83, c1_n21_w84, c1_n21_w85, c1_n21_w86, c1_n21_w87, c1_n21_w88, c1_n21_w89, c1_n21_w90, c1_n21_w91, c1_n21_w92, c1_n21_w93, c1_n21_w94, c1_n21_w95, c1_n21_w96, c1_n21_w97, c1_n21_w98, c1_n21_w99, c1_n21_w100, c1_n22_w1, c1_n22_w2, c1_n22_w3, c1_n22_w4, c1_n22_w5, c1_n22_w6, c1_n22_w7, c1_n22_w8, c1_n22_w9, c1_n22_w10, c1_n22_w11, c1_n22_w12, c1_n22_w13, c1_n22_w14, c1_n22_w15, c1_n22_w16, c1_n22_w17, c1_n22_w18, c1_n22_w19, c1_n22_w20, c1_n22_w21, c1_n22_w22, c1_n22_w23, c1_n22_w24, c1_n22_w25, c1_n22_w26, c1_n22_w27, c1_n22_w28, c1_n22_w29, c1_n22_w30, c1_n22_w31, c1_n22_w32, c1_n22_w33, c1_n22_w34, c1_n22_w35, c1_n22_w36, c1_n22_w37, c1_n22_w38, c1_n22_w39, c1_n22_w40, c1_n22_w41, c1_n22_w42, c1_n22_w43, c1_n22_w44, c1_n22_w45, c1_n22_w46, c1_n22_w47, c1_n22_w48, c1_n22_w49, c1_n22_w50, c1_n22_w51, c1_n22_w52, c1_n22_w53, c1_n22_w54, c1_n22_w55, c1_n22_w56, c1_n22_w57, c1_n22_w58, c1_n22_w59, c1_n22_w60, c1_n22_w61, c1_n22_w62, c1_n22_w63, c1_n22_w64, c1_n22_w65, c1_n22_w66, c1_n22_w67, c1_n22_w68, c1_n22_w69, c1_n22_w70, c1_n22_w71, c1_n22_w72, c1_n22_w73, c1_n22_w74, c1_n22_w75, c1_n22_w76, c1_n22_w77, c1_n22_w78, c1_n22_w79, c1_n22_w80, c1_n22_w81, c1_n22_w82, c1_n22_w83, c1_n22_w84, c1_n22_w85, c1_n22_w86, c1_n22_w87, c1_n22_w88, c1_n22_w89, c1_n22_w90, c1_n22_w91, c1_n22_w92, c1_n22_w93, c1_n22_w94, c1_n22_w95, c1_n22_w96, c1_n22_w97, c1_n22_w98, c1_n22_w99, c1_n22_w100, c1_n23_w1, c1_n23_w2, c1_n23_w3, c1_n23_w4, c1_n23_w5, c1_n23_w6, c1_n23_w7, c1_n23_w8, c1_n23_w9, c1_n23_w10, c1_n23_w11, c1_n23_w12, c1_n23_w13, c1_n23_w14, c1_n23_w15, c1_n23_w16, c1_n23_w17, c1_n23_w18, c1_n23_w19, c1_n23_w20, c1_n23_w21, c1_n23_w22, c1_n23_w23, c1_n23_w24, c1_n23_w25, c1_n23_w26, c1_n23_w27, c1_n23_w28, c1_n23_w29, c1_n23_w30, c1_n23_w31, c1_n23_w32, c1_n23_w33, c1_n23_w34, c1_n23_w35, c1_n23_w36, c1_n23_w37, c1_n23_w38, c1_n23_w39, c1_n23_w40, c1_n23_w41, c1_n23_w42, c1_n23_w43, c1_n23_w44, c1_n23_w45, c1_n23_w46, c1_n23_w47, c1_n23_w48, c1_n23_w49, c1_n23_w50, c1_n23_w51, c1_n23_w52, c1_n23_w53, c1_n23_w54, c1_n23_w55, c1_n23_w56, c1_n23_w57, c1_n23_w58, c1_n23_w59, c1_n23_w60, c1_n23_w61, c1_n23_w62, c1_n23_w63, c1_n23_w64, c1_n23_w65, c1_n23_w66, c1_n23_w67, c1_n23_w68, c1_n23_w69, c1_n23_w70, c1_n23_w71, c1_n23_w72, c1_n23_w73, c1_n23_w74, c1_n23_w75, c1_n23_w76, c1_n23_w77, c1_n23_w78, c1_n23_w79, c1_n23_w80, c1_n23_w81, c1_n23_w82, c1_n23_w83, c1_n23_w84, c1_n23_w85, c1_n23_w86, c1_n23_w87, c1_n23_w88, c1_n23_w89, c1_n23_w90, c1_n23_w91, c1_n23_w92, c1_n23_w93, c1_n23_w94, c1_n23_w95, c1_n23_w96, c1_n23_w97, c1_n23_w98, c1_n23_w99, c1_n23_w100, c1_n24_w1, c1_n24_w2, c1_n24_w3, c1_n24_w4, c1_n24_w5, c1_n24_w6, c1_n24_w7, c1_n24_w8, c1_n24_w9, c1_n24_w10, c1_n24_w11, c1_n24_w12, c1_n24_w13, c1_n24_w14, c1_n24_w15, c1_n24_w16, c1_n24_w17, c1_n24_w18, c1_n24_w19, c1_n24_w20, c1_n24_w21, c1_n24_w22, c1_n24_w23, c1_n24_w24, c1_n24_w25, c1_n24_w26, c1_n24_w27, c1_n24_w28, c1_n24_w29, c1_n24_w30, c1_n24_w31, c1_n24_w32, c1_n24_w33, c1_n24_w34, c1_n24_w35, c1_n24_w36, c1_n24_w37, c1_n24_w38, c1_n24_w39, c1_n24_w40, c1_n24_w41, c1_n24_w42, c1_n24_w43, c1_n24_w44, c1_n24_w45, c1_n24_w46, c1_n24_w47, c1_n24_w48, c1_n24_w49, c1_n24_w50, c1_n24_w51, c1_n24_w52, c1_n24_w53, c1_n24_w54, c1_n24_w55, c1_n24_w56, c1_n24_w57, c1_n24_w58, c1_n24_w59, c1_n24_w60, c1_n24_w61, c1_n24_w62, c1_n24_w63, c1_n24_w64, c1_n24_w65, c1_n24_w66, c1_n24_w67, c1_n24_w68, c1_n24_w69, c1_n24_w70, c1_n24_w71, c1_n24_w72, c1_n24_w73, c1_n24_w74, c1_n24_w75, c1_n24_w76, c1_n24_w77, c1_n24_w78, c1_n24_w79, c1_n24_w80, c1_n24_w81, c1_n24_w82, c1_n24_w83, c1_n24_w84, c1_n24_w85, c1_n24_w86, c1_n24_w87, c1_n24_w88, c1_n24_w89, c1_n24_w90, c1_n24_w91, c1_n24_w92, c1_n24_w93, c1_n24_w94, c1_n24_w95, c1_n24_w96, c1_n24_w97, c1_n24_w98, c1_n24_w99, c1_n24_w100, c1_n25_w1, c1_n25_w2, c1_n25_w3, c1_n25_w4, c1_n25_w5, c1_n25_w6, c1_n25_w7, c1_n25_w8, c1_n25_w9, c1_n25_w10, c1_n25_w11, c1_n25_w12, c1_n25_w13, c1_n25_w14, c1_n25_w15, c1_n25_w16, c1_n25_w17, c1_n25_w18, c1_n25_w19, c1_n25_w20, c1_n25_w21, c1_n25_w22, c1_n25_w23, c1_n25_w24, c1_n25_w25, c1_n25_w26, c1_n25_w27, c1_n25_w28, c1_n25_w29, c1_n25_w30, c1_n25_w31, c1_n25_w32, c1_n25_w33, c1_n25_w34, c1_n25_w35, c1_n25_w36, c1_n25_w37, c1_n25_w38, c1_n25_w39, c1_n25_w40, c1_n25_w41, c1_n25_w42, c1_n25_w43, c1_n25_w44, c1_n25_w45, c1_n25_w46, c1_n25_w47, c1_n25_w48, c1_n25_w49, c1_n25_w50, c1_n25_w51, c1_n25_w52, c1_n25_w53, c1_n25_w54, c1_n25_w55, c1_n25_w56, c1_n25_w57, c1_n25_w58, c1_n25_w59, c1_n25_w60, c1_n25_w61, c1_n25_w62, c1_n25_w63, c1_n25_w64, c1_n25_w65, c1_n25_w66, c1_n25_w67, c1_n25_w68, c1_n25_w69, c1_n25_w70, c1_n25_w71, c1_n25_w72, c1_n25_w73, c1_n25_w74, c1_n25_w75, c1_n25_w76, c1_n25_w77, c1_n25_w78, c1_n25_w79, c1_n25_w80, c1_n25_w81, c1_n25_w82, c1_n25_w83, c1_n25_w84, c1_n25_w85, c1_n25_w86, c1_n25_w87, c1_n25_w88, c1_n25_w89, c1_n25_w90, c1_n25_w91, c1_n25_w92, c1_n25_w93, c1_n25_w94, c1_n25_w95, c1_n25_w96, c1_n25_w97, c1_n25_w98, c1_n25_w99, c1_n25_w100, c1_n26_w1, c1_n26_w2, c1_n26_w3, c1_n26_w4, c1_n26_w5, c1_n26_w6, c1_n26_w7, c1_n26_w8, c1_n26_w9, c1_n26_w10, c1_n26_w11, c1_n26_w12, c1_n26_w13, c1_n26_w14, c1_n26_w15, c1_n26_w16, c1_n26_w17, c1_n26_w18, c1_n26_w19, c1_n26_w20, c1_n26_w21, c1_n26_w22, c1_n26_w23, c1_n26_w24, c1_n26_w25, c1_n26_w26, c1_n26_w27, c1_n26_w28, c1_n26_w29, c1_n26_w30, c1_n26_w31, c1_n26_w32, c1_n26_w33, c1_n26_w34, c1_n26_w35, c1_n26_w36, c1_n26_w37, c1_n26_w38, c1_n26_w39, c1_n26_w40, c1_n26_w41, c1_n26_w42, c1_n26_w43, c1_n26_w44, c1_n26_w45, c1_n26_w46, c1_n26_w47, c1_n26_w48, c1_n26_w49, c1_n26_w50, c1_n26_w51, c1_n26_w52, c1_n26_w53, c1_n26_w54, c1_n26_w55, c1_n26_w56, c1_n26_w57, c1_n26_w58, c1_n26_w59, c1_n26_w60, c1_n26_w61, c1_n26_w62, c1_n26_w63, c1_n26_w64, c1_n26_w65, c1_n26_w66, c1_n26_w67, c1_n26_w68, c1_n26_w69, c1_n26_w70, c1_n26_w71, c1_n26_w72, c1_n26_w73, c1_n26_w74, c1_n26_w75, c1_n26_w76, c1_n26_w77, c1_n26_w78, c1_n26_w79, c1_n26_w80, c1_n26_w81, c1_n26_w82, c1_n26_w83, c1_n26_w84, c1_n26_w85, c1_n26_w86, c1_n26_w87, c1_n26_w88, c1_n26_w89, c1_n26_w90, c1_n26_w91, c1_n26_w92, c1_n26_w93, c1_n26_w94, c1_n26_w95, c1_n26_w96, c1_n26_w97, c1_n26_w98, c1_n26_w99, c1_n26_w100, c1_n27_w1, c1_n27_w2, c1_n27_w3, c1_n27_w4, c1_n27_w5, c1_n27_w6, c1_n27_w7, c1_n27_w8, c1_n27_w9, c1_n27_w10, c1_n27_w11, c1_n27_w12, c1_n27_w13, c1_n27_w14, c1_n27_w15, c1_n27_w16, c1_n27_w17, c1_n27_w18, c1_n27_w19, c1_n27_w20, c1_n27_w21, c1_n27_w22, c1_n27_w23, c1_n27_w24, c1_n27_w25, c1_n27_w26, c1_n27_w27, c1_n27_w28, c1_n27_w29, c1_n27_w30, c1_n27_w31, c1_n27_w32, c1_n27_w33, c1_n27_w34, c1_n27_w35, c1_n27_w36, c1_n27_w37, c1_n27_w38, c1_n27_w39, c1_n27_w40, c1_n27_w41, c1_n27_w42, c1_n27_w43, c1_n27_w44, c1_n27_w45, c1_n27_w46, c1_n27_w47, c1_n27_w48, c1_n27_w49, c1_n27_w50, c1_n27_w51, c1_n27_w52, c1_n27_w53, c1_n27_w54, c1_n27_w55, c1_n27_w56, c1_n27_w57, c1_n27_w58, c1_n27_w59, c1_n27_w60, c1_n27_w61, c1_n27_w62, c1_n27_w63, c1_n27_w64, c1_n27_w65, c1_n27_w66, c1_n27_w67, c1_n27_w68, c1_n27_w69, c1_n27_w70, c1_n27_w71, c1_n27_w72, c1_n27_w73, c1_n27_w74, c1_n27_w75, c1_n27_w76, c1_n27_w77, c1_n27_w78, c1_n27_w79, c1_n27_w80, c1_n27_w81, c1_n27_w82, c1_n27_w83, c1_n27_w84, c1_n27_w85, c1_n27_w86, c1_n27_w87, c1_n27_w88, c1_n27_w89, c1_n27_w90, c1_n27_w91, c1_n27_w92, c1_n27_w93, c1_n27_w94, c1_n27_w95, c1_n27_w96, c1_n27_w97, c1_n27_w98, c1_n27_w99, c1_n27_w100, c1_n28_w1, c1_n28_w2, c1_n28_w3, c1_n28_w4, c1_n28_w5, c1_n28_w6, c1_n28_w7, c1_n28_w8, c1_n28_w9, c1_n28_w10, c1_n28_w11, c1_n28_w12, c1_n28_w13, c1_n28_w14, c1_n28_w15, c1_n28_w16, c1_n28_w17, c1_n28_w18, c1_n28_w19, c1_n28_w20, c1_n28_w21, c1_n28_w22, c1_n28_w23, c1_n28_w24, c1_n28_w25, c1_n28_w26, c1_n28_w27, c1_n28_w28, c1_n28_w29, c1_n28_w30, c1_n28_w31, c1_n28_w32, c1_n28_w33, c1_n28_w34, c1_n28_w35, c1_n28_w36, c1_n28_w37, c1_n28_w38, c1_n28_w39, c1_n28_w40, c1_n28_w41, c1_n28_w42, c1_n28_w43, c1_n28_w44, c1_n28_w45, c1_n28_w46, c1_n28_w47, c1_n28_w48, c1_n28_w49, c1_n28_w50, c1_n28_w51, c1_n28_w52, c1_n28_w53, c1_n28_w54, c1_n28_w55, c1_n28_w56, c1_n28_w57, c1_n28_w58, c1_n28_w59, c1_n28_w60, c1_n28_w61, c1_n28_w62, c1_n28_w63, c1_n28_w64, c1_n28_w65, c1_n28_w66, c1_n28_w67, c1_n28_w68, c1_n28_w69, c1_n28_w70, c1_n28_w71, c1_n28_w72, c1_n28_w73, c1_n28_w74, c1_n28_w75, c1_n28_w76, c1_n28_w77, c1_n28_w78, c1_n28_w79, c1_n28_w80, c1_n28_w81, c1_n28_w82, c1_n28_w83, c1_n28_w84, c1_n28_w85, c1_n28_w86, c1_n28_w87, c1_n28_w88, c1_n28_w89, c1_n28_w90, c1_n28_w91, c1_n28_w92, c1_n28_w93, c1_n28_w94, c1_n28_w95, c1_n28_w96, c1_n28_w97, c1_n28_w98, c1_n28_w99, c1_n28_w100, c1_n29_w1, c1_n29_w2, c1_n29_w3, c1_n29_w4, c1_n29_w5, c1_n29_w6, c1_n29_w7, c1_n29_w8, c1_n29_w9, c1_n29_w10, c1_n29_w11, c1_n29_w12, c1_n29_w13, c1_n29_w14, c1_n29_w15, c1_n29_w16, c1_n29_w17, c1_n29_w18, c1_n29_w19, c1_n29_w20, c1_n29_w21, c1_n29_w22, c1_n29_w23, c1_n29_w24, c1_n29_w25, c1_n29_w26, c1_n29_w27, c1_n29_w28, c1_n29_w29, c1_n29_w30, c1_n29_w31, c1_n29_w32, c1_n29_w33, c1_n29_w34, c1_n29_w35, c1_n29_w36, c1_n29_w37, c1_n29_w38, c1_n29_w39, c1_n29_w40, c1_n29_w41, c1_n29_w42, c1_n29_w43, c1_n29_w44, c1_n29_w45, c1_n29_w46, c1_n29_w47, c1_n29_w48, c1_n29_w49, c1_n29_w50, c1_n29_w51, c1_n29_w52, c1_n29_w53, c1_n29_w54, c1_n29_w55, c1_n29_w56, c1_n29_w57, c1_n29_w58, c1_n29_w59, c1_n29_w60, c1_n29_w61, c1_n29_w62, c1_n29_w63, c1_n29_w64, c1_n29_w65, c1_n29_w66, c1_n29_w67, c1_n29_w68, c1_n29_w69, c1_n29_w70, c1_n29_w71, c1_n29_w72, c1_n29_w73, c1_n29_w74, c1_n29_w75, c1_n29_w76, c1_n29_w77, c1_n29_w78, c1_n29_w79, c1_n29_w80, c1_n29_w81, c1_n29_w82, c1_n29_w83, c1_n29_w84, c1_n29_w85, c1_n29_w86, c1_n29_w87, c1_n29_w88, c1_n29_w89, c1_n29_w90, c1_n29_w91, c1_n29_w92, c1_n29_w93, c1_n29_w94, c1_n29_w95, c1_n29_w96, c1_n29_w97, c1_n29_w98, c1_n29_w99, c1_n29_w100, c1_n30_w1, c1_n30_w2, c1_n30_w3, c1_n30_w4, c1_n30_w5, c1_n30_w6, c1_n30_w7, c1_n30_w8, c1_n30_w9, c1_n30_w10, c1_n30_w11, c1_n30_w12, c1_n30_w13, c1_n30_w14, c1_n30_w15, c1_n30_w16, c1_n30_w17, c1_n30_w18, c1_n30_w19, c1_n30_w20, c1_n30_w21, c1_n30_w22, c1_n30_w23, c1_n30_w24, c1_n30_w25, c1_n30_w26, c1_n30_w27, c1_n30_w28, c1_n30_w29, c1_n30_w30, c1_n30_w31, c1_n30_w32, c1_n30_w33, c1_n30_w34, c1_n30_w35, c1_n30_w36, c1_n30_w37, c1_n30_w38, c1_n30_w39, c1_n30_w40, c1_n30_w41, c1_n30_w42, c1_n30_w43, c1_n30_w44, c1_n30_w45, c1_n30_w46, c1_n30_w47, c1_n30_w48, c1_n30_w49, c1_n30_w50, c1_n30_w51, c1_n30_w52, c1_n30_w53, c1_n30_w54, c1_n30_w55, c1_n30_w56, c1_n30_w57, c1_n30_w58, c1_n30_w59, c1_n30_w60, c1_n30_w61, c1_n30_w62, c1_n30_w63, c1_n30_w64, c1_n30_w65, c1_n30_w66, c1_n30_w67, c1_n30_w68, c1_n30_w69, c1_n30_w70, c1_n30_w71, c1_n30_w72, c1_n30_w73, c1_n30_w74, c1_n30_w75, c1_n30_w76, c1_n30_w77, c1_n30_w78, c1_n30_w79, c1_n30_w80, c1_n30_w81, c1_n30_w82, c1_n30_w83, c1_n30_w84, c1_n30_w85, c1_n30_w86, c1_n30_w87, c1_n30_w88, c1_n30_w89, c1_n30_w90, c1_n30_w91, c1_n30_w92, c1_n30_w93, c1_n30_w94, c1_n30_w95, c1_n30_w96, c1_n30_w97, c1_n30_w98, c1_n30_w99, c1_n30_w100, c1_n31_w1, c1_n31_w2, c1_n31_w3, c1_n31_w4, c1_n31_w5, c1_n31_w6, c1_n31_w7, c1_n31_w8, c1_n31_w9, c1_n31_w10, c1_n31_w11, c1_n31_w12, c1_n31_w13, c1_n31_w14, c1_n31_w15, c1_n31_w16, c1_n31_w17, c1_n31_w18, c1_n31_w19, c1_n31_w20, c1_n31_w21, c1_n31_w22, c1_n31_w23, c1_n31_w24, c1_n31_w25, c1_n31_w26, c1_n31_w27, c1_n31_w28, c1_n31_w29, c1_n31_w30, c1_n31_w31, c1_n31_w32, c1_n31_w33, c1_n31_w34, c1_n31_w35, c1_n31_w36, c1_n31_w37, c1_n31_w38, c1_n31_w39, c1_n31_w40, c1_n31_w41, c1_n31_w42, c1_n31_w43, c1_n31_w44, c1_n31_w45, c1_n31_w46, c1_n31_w47, c1_n31_w48, c1_n31_w49, c1_n31_w50, c1_n31_w51, c1_n31_w52, c1_n31_w53, c1_n31_w54, c1_n31_w55, c1_n31_w56, c1_n31_w57, c1_n31_w58, c1_n31_w59, c1_n31_w60, c1_n31_w61, c1_n31_w62, c1_n31_w63, c1_n31_w64, c1_n31_w65, c1_n31_w66, c1_n31_w67, c1_n31_w68, c1_n31_w69, c1_n31_w70, c1_n31_w71, c1_n31_w72, c1_n31_w73, c1_n31_w74, c1_n31_w75, c1_n31_w76, c1_n31_w77, c1_n31_w78, c1_n31_w79, c1_n31_w80, c1_n31_w81, c1_n31_w82, c1_n31_w83, c1_n31_w84, c1_n31_w85, c1_n31_w86, c1_n31_w87, c1_n31_w88, c1_n31_w89, c1_n31_w90, c1_n31_w91, c1_n31_w92, c1_n31_w93, c1_n31_w94, c1_n31_w95, c1_n31_w96, c1_n31_w97, c1_n31_w98, c1_n31_w99, c1_n31_w100, c1_n32_w1, c1_n32_w2, c1_n32_w3, c1_n32_w4, c1_n32_w5, c1_n32_w6, c1_n32_w7, c1_n32_w8, c1_n32_w9, c1_n32_w10, c1_n32_w11, c1_n32_w12, c1_n32_w13, c1_n32_w14, c1_n32_w15, c1_n32_w16, c1_n32_w17, c1_n32_w18, c1_n32_w19, c1_n32_w20, c1_n32_w21, c1_n32_w22, c1_n32_w23, c1_n32_w24, c1_n32_w25, c1_n32_w26, c1_n32_w27, c1_n32_w28, c1_n32_w29, c1_n32_w30, c1_n32_w31, c1_n32_w32, c1_n32_w33, c1_n32_w34, c1_n32_w35, c1_n32_w36, c1_n32_w37, c1_n32_w38, c1_n32_w39, c1_n32_w40, c1_n32_w41, c1_n32_w42, c1_n32_w43, c1_n32_w44, c1_n32_w45, c1_n32_w46, c1_n32_w47, c1_n32_w48, c1_n32_w49, c1_n32_w50, c1_n32_w51, c1_n32_w52, c1_n32_w53, c1_n32_w54, c1_n32_w55, c1_n32_w56, c1_n32_w57, c1_n32_w58, c1_n32_w59, c1_n32_w60, c1_n32_w61, c1_n32_w62, c1_n32_w63, c1_n32_w64, c1_n32_w65, c1_n32_w66, c1_n32_w67, c1_n32_w68, c1_n32_w69, c1_n32_w70, c1_n32_w71, c1_n32_w72, c1_n32_w73, c1_n32_w74, c1_n32_w75, c1_n32_w76, c1_n32_w77, c1_n32_w78, c1_n32_w79, c1_n32_w80, c1_n32_w81, c1_n32_w82, c1_n32_w83, c1_n32_w84, c1_n32_w85, c1_n32_w86, c1_n32_w87, c1_n32_w88, c1_n32_w89, c1_n32_w90, c1_n32_w91, c1_n32_w92, c1_n32_w93, c1_n32_w94, c1_n32_w95, c1_n32_w96, c1_n32_w97, c1_n32_w98, c1_n32_w99, c1_n32_w100, c1_n33_w1, c1_n33_w2, c1_n33_w3, c1_n33_w4, c1_n33_w5, c1_n33_w6, c1_n33_w7, c1_n33_w8, c1_n33_w9, c1_n33_w10, c1_n33_w11, c1_n33_w12, c1_n33_w13, c1_n33_w14, c1_n33_w15, c1_n33_w16, c1_n33_w17, c1_n33_w18, c1_n33_w19, c1_n33_w20, c1_n33_w21, c1_n33_w22, c1_n33_w23, c1_n33_w24, c1_n33_w25, c1_n33_w26, c1_n33_w27, c1_n33_w28, c1_n33_w29, c1_n33_w30, c1_n33_w31, c1_n33_w32, c1_n33_w33, c1_n33_w34, c1_n33_w35, c1_n33_w36, c1_n33_w37, c1_n33_w38, c1_n33_w39, c1_n33_w40, c1_n33_w41, c1_n33_w42, c1_n33_w43, c1_n33_w44, c1_n33_w45, c1_n33_w46, c1_n33_w47, c1_n33_w48, c1_n33_w49, c1_n33_w50, c1_n33_w51, c1_n33_w52, c1_n33_w53, c1_n33_w54, c1_n33_w55, c1_n33_w56, c1_n33_w57, c1_n33_w58, c1_n33_w59, c1_n33_w60, c1_n33_w61, c1_n33_w62, c1_n33_w63, c1_n33_w64, c1_n33_w65, c1_n33_w66, c1_n33_w67, c1_n33_w68, c1_n33_w69, c1_n33_w70, c1_n33_w71, c1_n33_w72, c1_n33_w73, c1_n33_w74, c1_n33_w75, c1_n33_w76, c1_n33_w77, c1_n33_w78, c1_n33_w79, c1_n33_w80, c1_n33_w81, c1_n33_w82, c1_n33_w83, c1_n33_w84, c1_n33_w85, c1_n33_w86, c1_n33_w87, c1_n33_w88, c1_n33_w89, c1_n33_w90, c1_n33_w91, c1_n33_w92, c1_n33_w93, c1_n33_w94, c1_n33_w95, c1_n33_w96, c1_n33_w97, c1_n33_w98, c1_n33_w99, c1_n33_w100, c1_n34_w1, c1_n34_w2, c1_n34_w3, c1_n34_w4, c1_n34_w5, c1_n34_w6, c1_n34_w7, c1_n34_w8, c1_n34_w9, c1_n34_w10, c1_n34_w11, c1_n34_w12, c1_n34_w13, c1_n34_w14, c1_n34_w15, c1_n34_w16, c1_n34_w17, c1_n34_w18, c1_n34_w19, c1_n34_w20, c1_n34_w21, c1_n34_w22, c1_n34_w23, c1_n34_w24, c1_n34_w25, c1_n34_w26, c1_n34_w27, c1_n34_w28, c1_n34_w29, c1_n34_w30, c1_n34_w31, c1_n34_w32, c1_n34_w33, c1_n34_w34, c1_n34_w35, c1_n34_w36, c1_n34_w37, c1_n34_w38, c1_n34_w39, c1_n34_w40, c1_n34_w41, c1_n34_w42, c1_n34_w43, c1_n34_w44, c1_n34_w45, c1_n34_w46, c1_n34_w47, c1_n34_w48, c1_n34_w49, c1_n34_w50, c1_n34_w51, c1_n34_w52, c1_n34_w53, c1_n34_w54, c1_n34_w55, c1_n34_w56, c1_n34_w57, c1_n34_w58, c1_n34_w59, c1_n34_w60, c1_n34_w61, c1_n34_w62, c1_n34_w63, c1_n34_w64, c1_n34_w65, c1_n34_w66, c1_n34_w67, c1_n34_w68, c1_n34_w69, c1_n34_w70, c1_n34_w71, c1_n34_w72, c1_n34_w73, c1_n34_w74, c1_n34_w75, c1_n34_w76, c1_n34_w77, c1_n34_w78, c1_n34_w79, c1_n34_w80, c1_n34_w81, c1_n34_w82, c1_n34_w83, c1_n34_w84, c1_n34_w85, c1_n34_w86, c1_n34_w87, c1_n34_w88, c1_n34_w89, c1_n34_w90, c1_n34_w91, c1_n34_w92, c1_n34_w93, c1_n34_w94, c1_n34_w95, c1_n34_w96, c1_n34_w97, c1_n34_w98, c1_n34_w99, c1_n34_w100, c1_n35_w1, c1_n35_w2, c1_n35_w3, c1_n35_w4, c1_n35_w5, c1_n35_w6, c1_n35_w7, c1_n35_w8, c1_n35_w9, c1_n35_w10, c1_n35_w11, c1_n35_w12, c1_n35_w13, c1_n35_w14, c1_n35_w15, c1_n35_w16, c1_n35_w17, c1_n35_w18, c1_n35_w19, c1_n35_w20, c1_n35_w21, c1_n35_w22, c1_n35_w23, c1_n35_w24, c1_n35_w25, c1_n35_w26, c1_n35_w27, c1_n35_w28, c1_n35_w29, c1_n35_w30, c1_n35_w31, c1_n35_w32, c1_n35_w33, c1_n35_w34, c1_n35_w35, c1_n35_w36, c1_n35_w37, c1_n35_w38, c1_n35_w39, c1_n35_w40, c1_n35_w41, c1_n35_w42, c1_n35_w43, c1_n35_w44, c1_n35_w45, c1_n35_w46, c1_n35_w47, c1_n35_w48, c1_n35_w49, c1_n35_w50, c1_n35_w51, c1_n35_w52, c1_n35_w53, c1_n35_w54, c1_n35_w55, c1_n35_w56, c1_n35_w57, c1_n35_w58, c1_n35_w59, c1_n35_w60, c1_n35_w61, c1_n35_w62, c1_n35_w63, c1_n35_w64, c1_n35_w65, c1_n35_w66, c1_n35_w67, c1_n35_w68, c1_n35_w69, c1_n35_w70, c1_n35_w71, c1_n35_w72, c1_n35_w73, c1_n35_w74, c1_n35_w75, c1_n35_w76, c1_n35_w77, c1_n35_w78, c1_n35_w79, c1_n35_w80, c1_n35_w81, c1_n35_w82, c1_n35_w83, c1_n35_w84, c1_n35_w85, c1_n35_w86, c1_n35_w87, c1_n35_w88, c1_n35_w89, c1_n35_w90, c1_n35_w91, c1_n35_w92, c1_n35_w93, c1_n35_w94, c1_n35_w95, c1_n35_w96, c1_n35_w97, c1_n35_w98, c1_n35_w99, c1_n35_w100, c1_n36_w1, c1_n36_w2, c1_n36_w3, c1_n36_w4, c1_n36_w5, c1_n36_w6, c1_n36_w7, c1_n36_w8, c1_n36_w9, c1_n36_w10, c1_n36_w11, c1_n36_w12, c1_n36_w13, c1_n36_w14, c1_n36_w15, c1_n36_w16, c1_n36_w17, c1_n36_w18, c1_n36_w19, c1_n36_w20, c1_n36_w21, c1_n36_w22, c1_n36_w23, c1_n36_w24, c1_n36_w25, c1_n36_w26, c1_n36_w27, c1_n36_w28, c1_n36_w29, c1_n36_w30, c1_n36_w31, c1_n36_w32, c1_n36_w33, c1_n36_w34, c1_n36_w35, c1_n36_w36, c1_n36_w37, c1_n36_w38, c1_n36_w39, c1_n36_w40, c1_n36_w41, c1_n36_w42, c1_n36_w43, c1_n36_w44, c1_n36_w45, c1_n36_w46, c1_n36_w47, c1_n36_w48, c1_n36_w49, c1_n36_w50, c1_n36_w51, c1_n36_w52, c1_n36_w53, c1_n36_w54, c1_n36_w55, c1_n36_w56, c1_n36_w57, c1_n36_w58, c1_n36_w59, c1_n36_w60, c1_n36_w61, c1_n36_w62, c1_n36_w63, c1_n36_w64, c1_n36_w65, c1_n36_w66, c1_n36_w67, c1_n36_w68, c1_n36_w69, c1_n36_w70, c1_n36_w71, c1_n36_w72, c1_n36_w73, c1_n36_w74, c1_n36_w75, c1_n36_w76, c1_n36_w77, c1_n36_w78, c1_n36_w79, c1_n36_w80, c1_n36_w81, c1_n36_w82, c1_n36_w83, c1_n36_w84, c1_n36_w85, c1_n36_w86, c1_n36_w87, c1_n36_w88, c1_n36_w89, c1_n36_w90, c1_n36_w91, c1_n36_w92, c1_n36_w93, c1_n36_w94, c1_n36_w95, c1_n36_w96, c1_n36_w97, c1_n36_w98, c1_n36_w99, c1_n36_w100, c1_n37_w1, c1_n37_w2, c1_n37_w3, c1_n37_w4, c1_n37_w5, c1_n37_w6, c1_n37_w7, c1_n37_w8, c1_n37_w9, c1_n37_w10, c1_n37_w11, c1_n37_w12, c1_n37_w13, c1_n37_w14, c1_n37_w15, c1_n37_w16, c1_n37_w17, c1_n37_w18, c1_n37_w19, c1_n37_w20, c1_n37_w21, c1_n37_w22, c1_n37_w23, c1_n37_w24, c1_n37_w25, c1_n37_w26, c1_n37_w27, c1_n37_w28, c1_n37_w29, c1_n37_w30, c1_n37_w31, c1_n37_w32, c1_n37_w33, c1_n37_w34, c1_n37_w35, c1_n37_w36, c1_n37_w37, c1_n37_w38, c1_n37_w39, c1_n37_w40, c1_n37_w41, c1_n37_w42, c1_n37_w43, c1_n37_w44, c1_n37_w45, c1_n37_w46, c1_n37_w47, c1_n37_w48, c1_n37_w49, c1_n37_w50, c1_n37_w51, c1_n37_w52, c1_n37_w53, c1_n37_w54, c1_n37_w55, c1_n37_w56, c1_n37_w57, c1_n37_w58, c1_n37_w59, c1_n37_w60, c1_n37_w61, c1_n37_w62, c1_n37_w63, c1_n37_w64, c1_n37_w65, c1_n37_w66, c1_n37_w67, c1_n37_w68, c1_n37_w69, c1_n37_w70, c1_n37_w71, c1_n37_w72, c1_n37_w73, c1_n37_w74, c1_n37_w75, c1_n37_w76, c1_n37_w77, c1_n37_w78, c1_n37_w79, c1_n37_w80, c1_n37_w81, c1_n37_w82, c1_n37_w83, c1_n37_w84, c1_n37_w85, c1_n37_w86, c1_n37_w87, c1_n37_w88, c1_n37_w89, c1_n37_w90, c1_n37_w91, c1_n37_w92, c1_n37_w93, c1_n37_w94, c1_n37_w95, c1_n37_w96, c1_n37_w97, c1_n37_w98, c1_n37_w99, c1_n37_w100, c1_n38_w1, c1_n38_w2, c1_n38_w3, c1_n38_w4, c1_n38_w5, c1_n38_w6, c1_n38_w7, c1_n38_w8, c1_n38_w9, c1_n38_w10, c1_n38_w11, c1_n38_w12, c1_n38_w13, c1_n38_w14, c1_n38_w15, c1_n38_w16, c1_n38_w17, c1_n38_w18, c1_n38_w19, c1_n38_w20, c1_n38_w21, c1_n38_w22, c1_n38_w23, c1_n38_w24, c1_n38_w25, c1_n38_w26, c1_n38_w27, c1_n38_w28, c1_n38_w29, c1_n38_w30, c1_n38_w31, c1_n38_w32, c1_n38_w33, c1_n38_w34, c1_n38_w35, c1_n38_w36, c1_n38_w37, c1_n38_w38, c1_n38_w39, c1_n38_w40, c1_n38_w41, c1_n38_w42, c1_n38_w43, c1_n38_w44, c1_n38_w45, c1_n38_w46, c1_n38_w47, c1_n38_w48, c1_n38_w49, c1_n38_w50, c1_n38_w51, c1_n38_w52, c1_n38_w53, c1_n38_w54, c1_n38_w55, c1_n38_w56, c1_n38_w57, c1_n38_w58, c1_n38_w59, c1_n38_w60, c1_n38_w61, c1_n38_w62, c1_n38_w63, c1_n38_w64, c1_n38_w65, c1_n38_w66, c1_n38_w67, c1_n38_w68, c1_n38_w69, c1_n38_w70, c1_n38_w71, c1_n38_w72, c1_n38_w73, c1_n38_w74, c1_n38_w75, c1_n38_w76, c1_n38_w77, c1_n38_w78, c1_n38_w79, c1_n38_w80, c1_n38_w81, c1_n38_w82, c1_n38_w83, c1_n38_w84, c1_n38_w85, c1_n38_w86, c1_n38_w87, c1_n38_w88, c1_n38_w89, c1_n38_w90, c1_n38_w91, c1_n38_w92, c1_n38_w93, c1_n38_w94, c1_n38_w95, c1_n38_w96, c1_n38_w97, c1_n38_w98, c1_n38_w99, c1_n38_w100, c1_n39_w1, c1_n39_w2, c1_n39_w3, c1_n39_w4, c1_n39_w5, c1_n39_w6, c1_n39_w7, c1_n39_w8, c1_n39_w9, c1_n39_w10, c1_n39_w11, c1_n39_w12, c1_n39_w13, c1_n39_w14, c1_n39_w15, c1_n39_w16, c1_n39_w17, c1_n39_w18, c1_n39_w19, c1_n39_w20, c1_n39_w21, c1_n39_w22, c1_n39_w23, c1_n39_w24, c1_n39_w25, c1_n39_w26, c1_n39_w27, c1_n39_w28, c1_n39_w29, c1_n39_w30, c1_n39_w31, c1_n39_w32, c1_n39_w33, c1_n39_w34, c1_n39_w35, c1_n39_w36, c1_n39_w37, c1_n39_w38, c1_n39_w39, c1_n39_w40, c1_n39_w41, c1_n39_w42, c1_n39_w43, c1_n39_w44, c1_n39_w45, c1_n39_w46, c1_n39_w47, c1_n39_w48, c1_n39_w49, c1_n39_w50, c1_n39_w51, c1_n39_w52, c1_n39_w53, c1_n39_w54, c1_n39_w55, c1_n39_w56, c1_n39_w57, c1_n39_w58, c1_n39_w59, c1_n39_w60, c1_n39_w61, c1_n39_w62, c1_n39_w63, c1_n39_w64, c1_n39_w65, c1_n39_w66, c1_n39_w67, c1_n39_w68, c1_n39_w69, c1_n39_w70, c1_n39_w71, c1_n39_w72, c1_n39_w73, c1_n39_w74, c1_n39_w75, c1_n39_w76, c1_n39_w77, c1_n39_w78, c1_n39_w79, c1_n39_w80, c1_n39_w81, c1_n39_w82, c1_n39_w83, c1_n39_w84, c1_n39_w85, c1_n39_w86, c1_n39_w87, c1_n39_w88, c1_n39_w89, c1_n39_w90, c1_n39_w91, c1_n39_w92, c1_n39_w93, c1_n39_w94, c1_n39_w95, c1_n39_w96, c1_n39_w97, c1_n39_w98, c1_n39_w99, c1_n39_w100, c1_n40_w1, c1_n40_w2, c1_n40_w3, c1_n40_w4, c1_n40_w5, c1_n40_w6, c1_n40_w7, c1_n40_w8, c1_n40_w9, c1_n40_w10, c1_n40_w11, c1_n40_w12, c1_n40_w13, c1_n40_w14, c1_n40_w15, c1_n40_w16, c1_n40_w17, c1_n40_w18, c1_n40_w19, c1_n40_w20, c1_n40_w21, c1_n40_w22, c1_n40_w23, c1_n40_w24, c1_n40_w25, c1_n40_w26, c1_n40_w27, c1_n40_w28, c1_n40_w29, c1_n40_w30, c1_n40_w31, c1_n40_w32, c1_n40_w33, c1_n40_w34, c1_n40_w35, c1_n40_w36, c1_n40_w37, c1_n40_w38, c1_n40_w39, c1_n40_w40, c1_n40_w41, c1_n40_w42, c1_n40_w43, c1_n40_w44, c1_n40_w45, c1_n40_w46, c1_n40_w47, c1_n40_w48, c1_n40_w49, c1_n40_w50, c1_n40_w51, c1_n40_w52, c1_n40_w53, c1_n40_w54, c1_n40_w55, c1_n40_w56, c1_n40_w57, c1_n40_w58, c1_n40_w59, c1_n40_w60, c1_n40_w61, c1_n40_w62, c1_n40_w63, c1_n40_w64, c1_n40_w65, c1_n40_w66, c1_n40_w67, c1_n40_w68, c1_n40_w69, c1_n40_w70, c1_n40_w71, c1_n40_w72, c1_n40_w73, c1_n40_w74, c1_n40_w75, c1_n40_w76, c1_n40_w77, c1_n40_w78, c1_n40_w79, c1_n40_w80, c1_n40_w81, c1_n40_w82, c1_n40_w83, c1_n40_w84, c1_n40_w85, c1_n40_w86, c1_n40_w87, c1_n40_w88, c1_n40_w89, c1_n40_w90, c1_n40_w91, c1_n40_w92, c1_n40_w93, c1_n40_w94, c1_n40_w95, c1_n40_w96, c1_n40_w97, c1_n40_w98, c1_n40_w99, c1_n40_w100, c1_n41_w1, c1_n41_w2, c1_n41_w3, c1_n41_w4, c1_n41_w5, c1_n41_w6, c1_n41_w7, c1_n41_w8, c1_n41_w9, c1_n41_w10, c1_n41_w11, c1_n41_w12, c1_n41_w13, c1_n41_w14, c1_n41_w15, c1_n41_w16, c1_n41_w17, c1_n41_w18, c1_n41_w19, c1_n41_w20, c1_n41_w21, c1_n41_w22, c1_n41_w23, c1_n41_w24, c1_n41_w25, c1_n41_w26, c1_n41_w27, c1_n41_w28, c1_n41_w29, c1_n41_w30, c1_n41_w31, c1_n41_w32, c1_n41_w33, c1_n41_w34, c1_n41_w35, c1_n41_w36, c1_n41_w37, c1_n41_w38, c1_n41_w39, c1_n41_w40, c1_n41_w41, c1_n41_w42, c1_n41_w43, c1_n41_w44, c1_n41_w45, c1_n41_w46, c1_n41_w47, c1_n41_w48, c1_n41_w49, c1_n41_w50, c1_n41_w51, c1_n41_w52, c1_n41_w53, c1_n41_w54, c1_n41_w55, c1_n41_w56, c1_n41_w57, c1_n41_w58, c1_n41_w59, c1_n41_w60, c1_n41_w61, c1_n41_w62, c1_n41_w63, c1_n41_w64, c1_n41_w65, c1_n41_w66, c1_n41_w67, c1_n41_w68, c1_n41_w69, c1_n41_w70, c1_n41_w71, c1_n41_w72, c1_n41_w73, c1_n41_w74, c1_n41_w75, c1_n41_w76, c1_n41_w77, c1_n41_w78, c1_n41_w79, c1_n41_w80, c1_n41_w81, c1_n41_w82, c1_n41_w83, c1_n41_w84, c1_n41_w85, c1_n41_w86, c1_n41_w87, c1_n41_w88, c1_n41_w89, c1_n41_w90, c1_n41_w91, c1_n41_w92, c1_n41_w93, c1_n41_w94, c1_n41_w95, c1_n41_w96, c1_n41_w97, c1_n41_w98, c1_n41_w99, c1_n41_w100, c1_n42_w1, c1_n42_w2, c1_n42_w3, c1_n42_w4, c1_n42_w5, c1_n42_w6, c1_n42_w7, c1_n42_w8, c1_n42_w9, c1_n42_w10, c1_n42_w11, c1_n42_w12, c1_n42_w13, c1_n42_w14, c1_n42_w15, c1_n42_w16, c1_n42_w17, c1_n42_w18, c1_n42_w19, c1_n42_w20, c1_n42_w21, c1_n42_w22, c1_n42_w23, c1_n42_w24, c1_n42_w25, c1_n42_w26, c1_n42_w27, c1_n42_w28, c1_n42_w29, c1_n42_w30, c1_n42_w31, c1_n42_w32, c1_n42_w33, c1_n42_w34, c1_n42_w35, c1_n42_w36, c1_n42_w37, c1_n42_w38, c1_n42_w39, c1_n42_w40, c1_n42_w41, c1_n42_w42, c1_n42_w43, c1_n42_w44, c1_n42_w45, c1_n42_w46, c1_n42_w47, c1_n42_w48, c1_n42_w49, c1_n42_w50, c1_n42_w51, c1_n42_w52, c1_n42_w53, c1_n42_w54, c1_n42_w55, c1_n42_w56, c1_n42_w57, c1_n42_w58, c1_n42_w59, c1_n42_w60, c1_n42_w61, c1_n42_w62, c1_n42_w63, c1_n42_w64, c1_n42_w65, c1_n42_w66, c1_n42_w67, c1_n42_w68, c1_n42_w69, c1_n42_w70, c1_n42_w71, c1_n42_w72, c1_n42_w73, c1_n42_w74, c1_n42_w75, c1_n42_w76, c1_n42_w77, c1_n42_w78, c1_n42_w79, c1_n42_w80, c1_n42_w81, c1_n42_w82, c1_n42_w83, c1_n42_w84, c1_n42_w85, c1_n42_w86, c1_n42_w87, c1_n42_w88, c1_n42_w89, c1_n42_w90, c1_n42_w91, c1_n42_w92, c1_n42_w93, c1_n42_w94, c1_n42_w95, c1_n42_w96, c1_n42_w97, c1_n42_w98, c1_n42_w99, c1_n42_w100, c1_n43_w1, c1_n43_w2, c1_n43_w3, c1_n43_w4, c1_n43_w5, c1_n43_w6, c1_n43_w7, c1_n43_w8, c1_n43_w9, c1_n43_w10, c1_n43_w11, c1_n43_w12, c1_n43_w13, c1_n43_w14, c1_n43_w15, c1_n43_w16, c1_n43_w17, c1_n43_w18, c1_n43_w19, c1_n43_w20, c1_n43_w21, c1_n43_w22, c1_n43_w23, c1_n43_w24, c1_n43_w25, c1_n43_w26, c1_n43_w27, c1_n43_w28, c1_n43_w29, c1_n43_w30, c1_n43_w31, c1_n43_w32, c1_n43_w33, c1_n43_w34, c1_n43_w35, c1_n43_w36, c1_n43_w37, c1_n43_w38, c1_n43_w39, c1_n43_w40, c1_n43_w41, c1_n43_w42, c1_n43_w43, c1_n43_w44, c1_n43_w45, c1_n43_w46, c1_n43_w47, c1_n43_w48, c1_n43_w49, c1_n43_w50, c1_n43_w51, c1_n43_w52, c1_n43_w53, c1_n43_w54, c1_n43_w55, c1_n43_w56, c1_n43_w57, c1_n43_w58, c1_n43_w59, c1_n43_w60, c1_n43_w61, c1_n43_w62, c1_n43_w63, c1_n43_w64, c1_n43_w65, c1_n43_w66, c1_n43_w67, c1_n43_w68, c1_n43_w69, c1_n43_w70, c1_n43_w71, c1_n43_w72, c1_n43_w73, c1_n43_w74, c1_n43_w75, c1_n43_w76, c1_n43_w77, c1_n43_w78, c1_n43_w79, c1_n43_w80, c1_n43_w81, c1_n43_w82, c1_n43_w83, c1_n43_w84, c1_n43_w85, c1_n43_w86, c1_n43_w87, c1_n43_w88, c1_n43_w89, c1_n43_w90, c1_n43_w91, c1_n43_w92, c1_n43_w93, c1_n43_w94, c1_n43_w95, c1_n43_w96, c1_n43_w97, c1_n43_w98, c1_n43_w99, c1_n43_w100, c1_n44_w1, c1_n44_w2, c1_n44_w3, c1_n44_w4, c1_n44_w5, c1_n44_w6, c1_n44_w7, c1_n44_w8, c1_n44_w9, c1_n44_w10, c1_n44_w11, c1_n44_w12, c1_n44_w13, c1_n44_w14, c1_n44_w15, c1_n44_w16, c1_n44_w17, c1_n44_w18, c1_n44_w19, c1_n44_w20, c1_n44_w21, c1_n44_w22, c1_n44_w23, c1_n44_w24, c1_n44_w25, c1_n44_w26, c1_n44_w27, c1_n44_w28, c1_n44_w29, c1_n44_w30, c1_n44_w31, c1_n44_w32, c1_n44_w33, c1_n44_w34, c1_n44_w35, c1_n44_w36, c1_n44_w37, c1_n44_w38, c1_n44_w39, c1_n44_w40, c1_n44_w41, c1_n44_w42, c1_n44_w43, c1_n44_w44, c1_n44_w45, c1_n44_w46, c1_n44_w47, c1_n44_w48, c1_n44_w49, c1_n44_w50, c1_n44_w51, c1_n44_w52, c1_n44_w53, c1_n44_w54, c1_n44_w55, c1_n44_w56, c1_n44_w57, c1_n44_w58, c1_n44_w59, c1_n44_w60, c1_n44_w61, c1_n44_w62, c1_n44_w63, c1_n44_w64, c1_n44_w65, c1_n44_w66, c1_n44_w67, c1_n44_w68, c1_n44_w69, c1_n44_w70, c1_n44_w71, c1_n44_w72, c1_n44_w73, c1_n44_w74, c1_n44_w75, c1_n44_w76, c1_n44_w77, c1_n44_w78, c1_n44_w79, c1_n44_w80, c1_n44_w81, c1_n44_w82, c1_n44_w83, c1_n44_w84, c1_n44_w85, c1_n44_w86, c1_n44_w87, c1_n44_w88, c1_n44_w89, c1_n44_w90, c1_n44_w91, c1_n44_w92, c1_n44_w93, c1_n44_w94, c1_n44_w95, c1_n44_w96, c1_n44_w97, c1_n44_w98, c1_n44_w99, c1_n44_w100, c1_n45_w1, c1_n45_w2, c1_n45_w3, c1_n45_w4, c1_n45_w5, c1_n45_w6, c1_n45_w7, c1_n45_w8, c1_n45_w9, c1_n45_w10, c1_n45_w11, c1_n45_w12, c1_n45_w13, c1_n45_w14, c1_n45_w15, c1_n45_w16, c1_n45_w17, c1_n45_w18, c1_n45_w19, c1_n45_w20, c1_n45_w21, c1_n45_w22, c1_n45_w23, c1_n45_w24, c1_n45_w25, c1_n45_w26, c1_n45_w27, c1_n45_w28, c1_n45_w29, c1_n45_w30, c1_n45_w31, c1_n45_w32, c1_n45_w33, c1_n45_w34, c1_n45_w35, c1_n45_w36, c1_n45_w37, c1_n45_w38, c1_n45_w39, c1_n45_w40, c1_n45_w41, c1_n45_w42, c1_n45_w43, c1_n45_w44, c1_n45_w45, c1_n45_w46, c1_n45_w47, c1_n45_w48, c1_n45_w49, c1_n45_w50, c1_n45_w51, c1_n45_w52, c1_n45_w53, c1_n45_w54, c1_n45_w55, c1_n45_w56, c1_n45_w57, c1_n45_w58, c1_n45_w59, c1_n45_w60, c1_n45_w61, c1_n45_w62, c1_n45_w63, c1_n45_w64, c1_n45_w65, c1_n45_w66, c1_n45_w67, c1_n45_w68, c1_n45_w69, c1_n45_w70, c1_n45_w71, c1_n45_w72, c1_n45_w73, c1_n45_w74, c1_n45_w75, c1_n45_w76, c1_n45_w77, c1_n45_w78, c1_n45_w79, c1_n45_w80, c1_n45_w81, c1_n45_w82, c1_n45_w83, c1_n45_w84, c1_n45_w85, c1_n45_w86, c1_n45_w87, c1_n45_w88, c1_n45_w89, c1_n45_w90, c1_n45_w91, c1_n45_w92, c1_n45_w93, c1_n45_w94, c1_n45_w95, c1_n45_w96, c1_n45_w97, c1_n45_w98, c1_n45_w99, c1_n45_w100, c1_n46_w1, c1_n46_w2, c1_n46_w3, c1_n46_w4, c1_n46_w5, c1_n46_w6, c1_n46_w7, c1_n46_w8, c1_n46_w9, c1_n46_w10, c1_n46_w11, c1_n46_w12, c1_n46_w13, c1_n46_w14, c1_n46_w15, c1_n46_w16, c1_n46_w17, c1_n46_w18, c1_n46_w19, c1_n46_w20, c1_n46_w21, c1_n46_w22, c1_n46_w23, c1_n46_w24, c1_n46_w25, c1_n46_w26, c1_n46_w27, c1_n46_w28, c1_n46_w29, c1_n46_w30, c1_n46_w31, c1_n46_w32, c1_n46_w33, c1_n46_w34, c1_n46_w35, c1_n46_w36, c1_n46_w37, c1_n46_w38, c1_n46_w39, c1_n46_w40, c1_n46_w41, c1_n46_w42, c1_n46_w43, c1_n46_w44, c1_n46_w45, c1_n46_w46, c1_n46_w47, c1_n46_w48, c1_n46_w49, c1_n46_w50, c1_n46_w51, c1_n46_w52, c1_n46_w53, c1_n46_w54, c1_n46_w55, c1_n46_w56, c1_n46_w57, c1_n46_w58, c1_n46_w59, c1_n46_w60, c1_n46_w61, c1_n46_w62, c1_n46_w63, c1_n46_w64, c1_n46_w65, c1_n46_w66, c1_n46_w67, c1_n46_w68, c1_n46_w69, c1_n46_w70, c1_n46_w71, c1_n46_w72, c1_n46_w73, c1_n46_w74, c1_n46_w75, c1_n46_w76, c1_n46_w77, c1_n46_w78, c1_n46_w79, c1_n46_w80, c1_n46_w81, c1_n46_w82, c1_n46_w83, c1_n46_w84, c1_n46_w85, c1_n46_w86, c1_n46_w87, c1_n46_w88, c1_n46_w89, c1_n46_w90, c1_n46_w91, c1_n46_w92, c1_n46_w93, c1_n46_w94, c1_n46_w95, c1_n46_w96, c1_n46_w97, c1_n46_w98, c1_n46_w99, c1_n46_w100, c1_n47_w1, c1_n47_w2, c1_n47_w3, c1_n47_w4, c1_n47_w5, c1_n47_w6, c1_n47_w7, c1_n47_w8, c1_n47_w9, c1_n47_w10, c1_n47_w11, c1_n47_w12, c1_n47_w13, c1_n47_w14, c1_n47_w15, c1_n47_w16, c1_n47_w17, c1_n47_w18, c1_n47_w19, c1_n47_w20, c1_n47_w21, c1_n47_w22, c1_n47_w23, c1_n47_w24, c1_n47_w25, c1_n47_w26, c1_n47_w27, c1_n47_w28, c1_n47_w29, c1_n47_w30, c1_n47_w31, c1_n47_w32, c1_n47_w33, c1_n47_w34, c1_n47_w35, c1_n47_w36, c1_n47_w37, c1_n47_w38, c1_n47_w39, c1_n47_w40, c1_n47_w41, c1_n47_w42, c1_n47_w43, c1_n47_w44, c1_n47_w45, c1_n47_w46, c1_n47_w47, c1_n47_w48, c1_n47_w49, c1_n47_w50, c1_n47_w51, c1_n47_w52, c1_n47_w53, c1_n47_w54, c1_n47_w55, c1_n47_w56, c1_n47_w57, c1_n47_w58, c1_n47_w59, c1_n47_w60, c1_n47_w61, c1_n47_w62, c1_n47_w63, c1_n47_w64, c1_n47_w65, c1_n47_w66, c1_n47_w67, c1_n47_w68, c1_n47_w69, c1_n47_w70, c1_n47_w71, c1_n47_w72, c1_n47_w73, c1_n47_w74, c1_n47_w75, c1_n47_w76, c1_n47_w77, c1_n47_w78, c1_n47_w79, c1_n47_w80, c1_n47_w81, c1_n47_w82, c1_n47_w83, c1_n47_w84, c1_n47_w85, c1_n47_w86, c1_n47_w87, c1_n47_w88, c1_n47_w89, c1_n47_w90, c1_n47_w91, c1_n47_w92, c1_n47_w93, c1_n47_w94, c1_n47_w95, c1_n47_w96, c1_n47_w97, c1_n47_w98, c1_n47_w99, c1_n47_w100, c1_n48_w1, c1_n48_w2, c1_n48_w3, c1_n48_w4, c1_n48_w5, c1_n48_w6, c1_n48_w7, c1_n48_w8, c1_n48_w9, c1_n48_w10, c1_n48_w11, c1_n48_w12, c1_n48_w13, c1_n48_w14, c1_n48_w15, c1_n48_w16, c1_n48_w17, c1_n48_w18, c1_n48_w19, c1_n48_w20, c1_n48_w21, c1_n48_w22, c1_n48_w23, c1_n48_w24, c1_n48_w25, c1_n48_w26, c1_n48_w27, c1_n48_w28, c1_n48_w29, c1_n48_w30, c1_n48_w31, c1_n48_w32, c1_n48_w33, c1_n48_w34, c1_n48_w35, c1_n48_w36, c1_n48_w37, c1_n48_w38, c1_n48_w39, c1_n48_w40, c1_n48_w41, c1_n48_w42, c1_n48_w43, c1_n48_w44, c1_n48_w45, c1_n48_w46, c1_n48_w47, c1_n48_w48, c1_n48_w49, c1_n48_w50, c1_n48_w51, c1_n48_w52, c1_n48_w53, c1_n48_w54, c1_n48_w55, c1_n48_w56, c1_n48_w57, c1_n48_w58, c1_n48_w59, c1_n48_w60, c1_n48_w61, c1_n48_w62, c1_n48_w63, c1_n48_w64, c1_n48_w65, c1_n48_w66, c1_n48_w67, c1_n48_w68, c1_n48_w69, c1_n48_w70, c1_n48_w71, c1_n48_w72, c1_n48_w73, c1_n48_w74, c1_n48_w75, c1_n48_w76, c1_n48_w77, c1_n48_w78, c1_n48_w79, c1_n48_w80, c1_n48_w81, c1_n48_w82, c1_n48_w83, c1_n48_w84, c1_n48_w85, c1_n48_w86, c1_n48_w87, c1_n48_w88, c1_n48_w89, c1_n48_w90, c1_n48_w91, c1_n48_w92, c1_n48_w93, c1_n48_w94, c1_n48_w95, c1_n48_w96, c1_n48_w97, c1_n48_w98, c1_n48_w99, c1_n48_w100, c1_n49_w1, c1_n49_w2, c1_n49_w3, c1_n49_w4, c1_n49_w5, c1_n49_w6, c1_n49_w7, c1_n49_w8, c1_n49_w9, c1_n49_w10, c1_n49_w11, c1_n49_w12, c1_n49_w13, c1_n49_w14, c1_n49_w15, c1_n49_w16, c1_n49_w17, c1_n49_w18, c1_n49_w19, c1_n49_w20, c1_n49_w21, c1_n49_w22, c1_n49_w23, c1_n49_w24, c1_n49_w25, c1_n49_w26, c1_n49_w27, c1_n49_w28, c1_n49_w29, c1_n49_w30, c1_n49_w31, c1_n49_w32, c1_n49_w33, c1_n49_w34, c1_n49_w35, c1_n49_w36, c1_n49_w37, c1_n49_w38, c1_n49_w39, c1_n49_w40, c1_n49_w41, c1_n49_w42, c1_n49_w43, c1_n49_w44, c1_n49_w45, c1_n49_w46, c1_n49_w47, c1_n49_w48, c1_n49_w49, c1_n49_w50, c1_n49_w51, c1_n49_w52, c1_n49_w53, c1_n49_w54, c1_n49_w55, c1_n49_w56, c1_n49_w57, c1_n49_w58, c1_n49_w59, c1_n49_w60, c1_n49_w61, c1_n49_w62, c1_n49_w63, c1_n49_w64, c1_n49_w65, c1_n49_w66, c1_n49_w67, c1_n49_w68, c1_n49_w69, c1_n49_w70, c1_n49_w71, c1_n49_w72, c1_n49_w73, c1_n49_w74, c1_n49_w75, c1_n49_w76, c1_n49_w77, c1_n49_w78, c1_n49_w79, c1_n49_w80, c1_n49_w81, c1_n49_w82, c1_n49_w83, c1_n49_w84, c1_n49_w85, c1_n49_w86, c1_n49_w87, c1_n49_w88, c1_n49_w89, c1_n49_w90, c1_n49_w91, c1_n49_w92, c1_n49_w93, c1_n49_w94, c1_n49_w95, c1_n49_w96, c1_n49_w97, c1_n49_w98, c1_n49_w99, c1_n49_w100: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c1_n0_y, c1_n1_y, c1_n2_y, c1_n3_y, c1_n4_y, c1_n5_y, c1_n6_y, c1_n7_y, c1_n8_y, c1_n9_y, c1_n10_y, c1_n11_y, c1_n12_y, c1_n13_y, c1_n14_y, c1_n15_y, c1_n16_y, c1_n17_y, c1_n18_y, c1_n19_y, c1_n20_y, c1_n21_y, c1_n22_y, c1_n23_y, c1_n24_y, c1_n25_y, c1_n26_y, c1_n27_y, c1_n28_y, c1_n29_y, c1_n30_y, c1_n31_y, c1_n32_y, c1_n33_y, c1_n34_y, c1_n35_y, c1_n36_y, c1_n37_y, c1_n38_y, c1_n39_y, c1_n40_y, c1_n41_y, c1_n42_y, c1_n43_y, c1_n44_y, c1_n45_y, c1_n46_y, c1_n47_y, c1_n48_y, c1_n49_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada1_ReLU_50neuron_8bits_100n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n0_w1, 
            w2=> c1_n0_w2, 
            w3=> c1_n0_w3, 
            w4=> c1_n0_w4, 
            w5=> c1_n0_w5, 
            w6=> c1_n0_w6, 
            w7=> c1_n0_w7, 
            w8=> c1_n0_w8, 
            w9=> c1_n0_w9, 
            w10=> c1_n0_w10, 
            w11=> c1_n0_w11, 
            w12=> c1_n0_w12, 
            w13=> c1_n0_w13, 
            w14=> c1_n0_w14, 
            w15=> c1_n0_w15, 
            w16=> c1_n0_w16, 
            w17=> c1_n0_w17, 
            w18=> c1_n0_w18, 
            w19=> c1_n0_w19, 
            w20=> c1_n0_w20, 
            w21=> c1_n0_w21, 
            w22=> c1_n0_w22, 
            w23=> c1_n0_w23, 
            w24=> c1_n0_w24, 
            w25=> c1_n0_w25, 
            w26=> c1_n0_w26, 
            w27=> c1_n0_w27, 
            w28=> c1_n0_w28, 
            w29=> c1_n0_w29, 
            w30=> c1_n0_w30, 
            w31=> c1_n0_w31, 
            w32=> c1_n0_w32, 
            w33=> c1_n0_w33, 
            w34=> c1_n0_w34, 
            w35=> c1_n0_w35, 
            w36=> c1_n0_w36, 
            w37=> c1_n0_w37, 
            w38=> c1_n0_w38, 
            w39=> c1_n0_w39, 
            w40=> c1_n0_w40, 
            w41=> c1_n0_w41, 
            w42=> c1_n0_w42, 
            w43=> c1_n0_w43, 
            w44=> c1_n0_w44, 
            w45=> c1_n0_w45, 
            w46=> c1_n0_w46, 
            w47=> c1_n0_w47, 
            w48=> c1_n0_w48, 
            w49=> c1_n0_w49, 
            w50=> c1_n0_w50, 
            w51=> c1_n0_w51, 
            w52=> c1_n0_w52, 
            w53=> c1_n0_w53, 
            w54=> c1_n0_w54, 
            w55=> c1_n0_w55, 
            w56=> c1_n0_w56, 
            w57=> c1_n0_w57, 
            w58=> c1_n0_w58, 
            w59=> c1_n0_w59, 
            w60=> c1_n0_w60, 
            w61=> c1_n0_w61, 
            w62=> c1_n0_w62, 
            w63=> c1_n0_w63, 
            w64=> c1_n0_w64, 
            w65=> c1_n0_w65, 
            w66=> c1_n0_w66, 
            w67=> c1_n0_w67, 
            w68=> c1_n0_w68, 
            w69=> c1_n0_w69, 
            w70=> c1_n0_w70, 
            w71=> c1_n0_w71, 
            w72=> c1_n0_w72, 
            w73=> c1_n0_w73, 
            w74=> c1_n0_w74, 
            w75=> c1_n0_w75, 
            w76=> c1_n0_w76, 
            w77=> c1_n0_w77, 
            w78=> c1_n0_w78, 
            w79=> c1_n0_w79, 
            w80=> c1_n0_w80, 
            w81=> c1_n0_w81, 
            w82=> c1_n0_w82, 
            w83=> c1_n0_w83, 
            w84=> c1_n0_w84, 
            w85=> c1_n0_w85, 
            w86=> c1_n0_w86, 
            w87=> c1_n0_w87, 
            w88=> c1_n0_w88, 
            w89=> c1_n0_w89, 
            w90=> c1_n0_w90, 
            w91=> c1_n0_w91, 
            w92=> c1_n0_w92, 
            w93=> c1_n0_w93, 
            w94=> c1_n0_w94, 
            w95=> c1_n0_w95, 
            w96=> c1_n0_w96, 
            w97=> c1_n0_w97, 
            w98=> c1_n0_w98, 
            w99=> c1_n0_w99, 
            w100=> c1_n0_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n1_w1, 
            w2=> c1_n1_w2, 
            w3=> c1_n1_w3, 
            w4=> c1_n1_w4, 
            w5=> c1_n1_w5, 
            w6=> c1_n1_w6, 
            w7=> c1_n1_w7, 
            w8=> c1_n1_w8, 
            w9=> c1_n1_w9, 
            w10=> c1_n1_w10, 
            w11=> c1_n1_w11, 
            w12=> c1_n1_w12, 
            w13=> c1_n1_w13, 
            w14=> c1_n1_w14, 
            w15=> c1_n1_w15, 
            w16=> c1_n1_w16, 
            w17=> c1_n1_w17, 
            w18=> c1_n1_w18, 
            w19=> c1_n1_w19, 
            w20=> c1_n1_w20, 
            w21=> c1_n1_w21, 
            w22=> c1_n1_w22, 
            w23=> c1_n1_w23, 
            w24=> c1_n1_w24, 
            w25=> c1_n1_w25, 
            w26=> c1_n1_w26, 
            w27=> c1_n1_w27, 
            w28=> c1_n1_w28, 
            w29=> c1_n1_w29, 
            w30=> c1_n1_w30, 
            w31=> c1_n1_w31, 
            w32=> c1_n1_w32, 
            w33=> c1_n1_w33, 
            w34=> c1_n1_w34, 
            w35=> c1_n1_w35, 
            w36=> c1_n1_w36, 
            w37=> c1_n1_w37, 
            w38=> c1_n1_w38, 
            w39=> c1_n1_w39, 
            w40=> c1_n1_w40, 
            w41=> c1_n1_w41, 
            w42=> c1_n1_w42, 
            w43=> c1_n1_w43, 
            w44=> c1_n1_w44, 
            w45=> c1_n1_w45, 
            w46=> c1_n1_w46, 
            w47=> c1_n1_w47, 
            w48=> c1_n1_w48, 
            w49=> c1_n1_w49, 
            w50=> c1_n1_w50, 
            w51=> c1_n1_w51, 
            w52=> c1_n1_w52, 
            w53=> c1_n1_w53, 
            w54=> c1_n1_w54, 
            w55=> c1_n1_w55, 
            w56=> c1_n1_w56, 
            w57=> c1_n1_w57, 
            w58=> c1_n1_w58, 
            w59=> c1_n1_w59, 
            w60=> c1_n1_w60, 
            w61=> c1_n1_w61, 
            w62=> c1_n1_w62, 
            w63=> c1_n1_w63, 
            w64=> c1_n1_w64, 
            w65=> c1_n1_w65, 
            w66=> c1_n1_w66, 
            w67=> c1_n1_w67, 
            w68=> c1_n1_w68, 
            w69=> c1_n1_w69, 
            w70=> c1_n1_w70, 
            w71=> c1_n1_w71, 
            w72=> c1_n1_w72, 
            w73=> c1_n1_w73, 
            w74=> c1_n1_w74, 
            w75=> c1_n1_w75, 
            w76=> c1_n1_w76, 
            w77=> c1_n1_w77, 
            w78=> c1_n1_w78, 
            w79=> c1_n1_w79, 
            w80=> c1_n1_w80, 
            w81=> c1_n1_w81, 
            w82=> c1_n1_w82, 
            w83=> c1_n1_w83, 
            w84=> c1_n1_w84, 
            w85=> c1_n1_w85, 
            w86=> c1_n1_w86, 
            w87=> c1_n1_w87, 
            w88=> c1_n1_w88, 
            w89=> c1_n1_w89, 
            w90=> c1_n1_w90, 
            w91=> c1_n1_w91, 
            w92=> c1_n1_w92, 
            w93=> c1_n1_w93, 
            w94=> c1_n1_w94, 
            w95=> c1_n1_w95, 
            w96=> c1_n1_w96, 
            w97=> c1_n1_w97, 
            w98=> c1_n1_w98, 
            w99=> c1_n1_w99, 
            w100=> c1_n1_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n2_w1, 
            w2=> c1_n2_w2, 
            w3=> c1_n2_w3, 
            w4=> c1_n2_w4, 
            w5=> c1_n2_w5, 
            w6=> c1_n2_w6, 
            w7=> c1_n2_w7, 
            w8=> c1_n2_w8, 
            w9=> c1_n2_w9, 
            w10=> c1_n2_w10, 
            w11=> c1_n2_w11, 
            w12=> c1_n2_w12, 
            w13=> c1_n2_w13, 
            w14=> c1_n2_w14, 
            w15=> c1_n2_w15, 
            w16=> c1_n2_w16, 
            w17=> c1_n2_w17, 
            w18=> c1_n2_w18, 
            w19=> c1_n2_w19, 
            w20=> c1_n2_w20, 
            w21=> c1_n2_w21, 
            w22=> c1_n2_w22, 
            w23=> c1_n2_w23, 
            w24=> c1_n2_w24, 
            w25=> c1_n2_w25, 
            w26=> c1_n2_w26, 
            w27=> c1_n2_w27, 
            w28=> c1_n2_w28, 
            w29=> c1_n2_w29, 
            w30=> c1_n2_w30, 
            w31=> c1_n2_w31, 
            w32=> c1_n2_w32, 
            w33=> c1_n2_w33, 
            w34=> c1_n2_w34, 
            w35=> c1_n2_w35, 
            w36=> c1_n2_w36, 
            w37=> c1_n2_w37, 
            w38=> c1_n2_w38, 
            w39=> c1_n2_w39, 
            w40=> c1_n2_w40, 
            w41=> c1_n2_w41, 
            w42=> c1_n2_w42, 
            w43=> c1_n2_w43, 
            w44=> c1_n2_w44, 
            w45=> c1_n2_w45, 
            w46=> c1_n2_w46, 
            w47=> c1_n2_w47, 
            w48=> c1_n2_w48, 
            w49=> c1_n2_w49, 
            w50=> c1_n2_w50, 
            w51=> c1_n2_w51, 
            w52=> c1_n2_w52, 
            w53=> c1_n2_w53, 
            w54=> c1_n2_w54, 
            w55=> c1_n2_w55, 
            w56=> c1_n2_w56, 
            w57=> c1_n2_w57, 
            w58=> c1_n2_w58, 
            w59=> c1_n2_w59, 
            w60=> c1_n2_w60, 
            w61=> c1_n2_w61, 
            w62=> c1_n2_w62, 
            w63=> c1_n2_w63, 
            w64=> c1_n2_w64, 
            w65=> c1_n2_w65, 
            w66=> c1_n2_w66, 
            w67=> c1_n2_w67, 
            w68=> c1_n2_w68, 
            w69=> c1_n2_w69, 
            w70=> c1_n2_w70, 
            w71=> c1_n2_w71, 
            w72=> c1_n2_w72, 
            w73=> c1_n2_w73, 
            w74=> c1_n2_w74, 
            w75=> c1_n2_w75, 
            w76=> c1_n2_w76, 
            w77=> c1_n2_w77, 
            w78=> c1_n2_w78, 
            w79=> c1_n2_w79, 
            w80=> c1_n2_w80, 
            w81=> c1_n2_w81, 
            w82=> c1_n2_w82, 
            w83=> c1_n2_w83, 
            w84=> c1_n2_w84, 
            w85=> c1_n2_w85, 
            w86=> c1_n2_w86, 
            w87=> c1_n2_w87, 
            w88=> c1_n2_w88, 
            w89=> c1_n2_w89, 
            w90=> c1_n2_w90, 
            w91=> c1_n2_w91, 
            w92=> c1_n2_w92, 
            w93=> c1_n2_w93, 
            w94=> c1_n2_w94, 
            w95=> c1_n2_w95, 
            w96=> c1_n2_w96, 
            w97=> c1_n2_w97, 
            w98=> c1_n2_w98, 
            w99=> c1_n2_w99, 
            w100=> c1_n2_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n3_w1, 
            w2=> c1_n3_w2, 
            w3=> c1_n3_w3, 
            w4=> c1_n3_w4, 
            w5=> c1_n3_w5, 
            w6=> c1_n3_w6, 
            w7=> c1_n3_w7, 
            w8=> c1_n3_w8, 
            w9=> c1_n3_w9, 
            w10=> c1_n3_w10, 
            w11=> c1_n3_w11, 
            w12=> c1_n3_w12, 
            w13=> c1_n3_w13, 
            w14=> c1_n3_w14, 
            w15=> c1_n3_w15, 
            w16=> c1_n3_w16, 
            w17=> c1_n3_w17, 
            w18=> c1_n3_w18, 
            w19=> c1_n3_w19, 
            w20=> c1_n3_w20, 
            w21=> c1_n3_w21, 
            w22=> c1_n3_w22, 
            w23=> c1_n3_w23, 
            w24=> c1_n3_w24, 
            w25=> c1_n3_w25, 
            w26=> c1_n3_w26, 
            w27=> c1_n3_w27, 
            w28=> c1_n3_w28, 
            w29=> c1_n3_w29, 
            w30=> c1_n3_w30, 
            w31=> c1_n3_w31, 
            w32=> c1_n3_w32, 
            w33=> c1_n3_w33, 
            w34=> c1_n3_w34, 
            w35=> c1_n3_w35, 
            w36=> c1_n3_w36, 
            w37=> c1_n3_w37, 
            w38=> c1_n3_w38, 
            w39=> c1_n3_w39, 
            w40=> c1_n3_w40, 
            w41=> c1_n3_w41, 
            w42=> c1_n3_w42, 
            w43=> c1_n3_w43, 
            w44=> c1_n3_w44, 
            w45=> c1_n3_w45, 
            w46=> c1_n3_w46, 
            w47=> c1_n3_w47, 
            w48=> c1_n3_w48, 
            w49=> c1_n3_w49, 
            w50=> c1_n3_w50, 
            w51=> c1_n3_w51, 
            w52=> c1_n3_w52, 
            w53=> c1_n3_w53, 
            w54=> c1_n3_w54, 
            w55=> c1_n3_w55, 
            w56=> c1_n3_w56, 
            w57=> c1_n3_w57, 
            w58=> c1_n3_w58, 
            w59=> c1_n3_w59, 
            w60=> c1_n3_w60, 
            w61=> c1_n3_w61, 
            w62=> c1_n3_w62, 
            w63=> c1_n3_w63, 
            w64=> c1_n3_w64, 
            w65=> c1_n3_w65, 
            w66=> c1_n3_w66, 
            w67=> c1_n3_w67, 
            w68=> c1_n3_w68, 
            w69=> c1_n3_w69, 
            w70=> c1_n3_w70, 
            w71=> c1_n3_w71, 
            w72=> c1_n3_w72, 
            w73=> c1_n3_w73, 
            w74=> c1_n3_w74, 
            w75=> c1_n3_w75, 
            w76=> c1_n3_w76, 
            w77=> c1_n3_w77, 
            w78=> c1_n3_w78, 
            w79=> c1_n3_w79, 
            w80=> c1_n3_w80, 
            w81=> c1_n3_w81, 
            w82=> c1_n3_w82, 
            w83=> c1_n3_w83, 
            w84=> c1_n3_w84, 
            w85=> c1_n3_w85, 
            w86=> c1_n3_w86, 
            w87=> c1_n3_w87, 
            w88=> c1_n3_w88, 
            w89=> c1_n3_w89, 
            w90=> c1_n3_w90, 
            w91=> c1_n3_w91, 
            w92=> c1_n3_w92, 
            w93=> c1_n3_w93, 
            w94=> c1_n3_w94, 
            w95=> c1_n3_w95, 
            w96=> c1_n3_w96, 
            w97=> c1_n3_w97, 
            w98=> c1_n3_w98, 
            w99=> c1_n3_w99, 
            w100=> c1_n3_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n4_w1, 
            w2=> c1_n4_w2, 
            w3=> c1_n4_w3, 
            w4=> c1_n4_w4, 
            w5=> c1_n4_w5, 
            w6=> c1_n4_w6, 
            w7=> c1_n4_w7, 
            w8=> c1_n4_w8, 
            w9=> c1_n4_w9, 
            w10=> c1_n4_w10, 
            w11=> c1_n4_w11, 
            w12=> c1_n4_w12, 
            w13=> c1_n4_w13, 
            w14=> c1_n4_w14, 
            w15=> c1_n4_w15, 
            w16=> c1_n4_w16, 
            w17=> c1_n4_w17, 
            w18=> c1_n4_w18, 
            w19=> c1_n4_w19, 
            w20=> c1_n4_w20, 
            w21=> c1_n4_w21, 
            w22=> c1_n4_w22, 
            w23=> c1_n4_w23, 
            w24=> c1_n4_w24, 
            w25=> c1_n4_w25, 
            w26=> c1_n4_w26, 
            w27=> c1_n4_w27, 
            w28=> c1_n4_w28, 
            w29=> c1_n4_w29, 
            w30=> c1_n4_w30, 
            w31=> c1_n4_w31, 
            w32=> c1_n4_w32, 
            w33=> c1_n4_w33, 
            w34=> c1_n4_w34, 
            w35=> c1_n4_w35, 
            w36=> c1_n4_w36, 
            w37=> c1_n4_w37, 
            w38=> c1_n4_w38, 
            w39=> c1_n4_w39, 
            w40=> c1_n4_w40, 
            w41=> c1_n4_w41, 
            w42=> c1_n4_w42, 
            w43=> c1_n4_w43, 
            w44=> c1_n4_w44, 
            w45=> c1_n4_w45, 
            w46=> c1_n4_w46, 
            w47=> c1_n4_w47, 
            w48=> c1_n4_w48, 
            w49=> c1_n4_w49, 
            w50=> c1_n4_w50, 
            w51=> c1_n4_w51, 
            w52=> c1_n4_w52, 
            w53=> c1_n4_w53, 
            w54=> c1_n4_w54, 
            w55=> c1_n4_w55, 
            w56=> c1_n4_w56, 
            w57=> c1_n4_w57, 
            w58=> c1_n4_w58, 
            w59=> c1_n4_w59, 
            w60=> c1_n4_w60, 
            w61=> c1_n4_w61, 
            w62=> c1_n4_w62, 
            w63=> c1_n4_w63, 
            w64=> c1_n4_w64, 
            w65=> c1_n4_w65, 
            w66=> c1_n4_w66, 
            w67=> c1_n4_w67, 
            w68=> c1_n4_w68, 
            w69=> c1_n4_w69, 
            w70=> c1_n4_w70, 
            w71=> c1_n4_w71, 
            w72=> c1_n4_w72, 
            w73=> c1_n4_w73, 
            w74=> c1_n4_w74, 
            w75=> c1_n4_w75, 
            w76=> c1_n4_w76, 
            w77=> c1_n4_w77, 
            w78=> c1_n4_w78, 
            w79=> c1_n4_w79, 
            w80=> c1_n4_w80, 
            w81=> c1_n4_w81, 
            w82=> c1_n4_w82, 
            w83=> c1_n4_w83, 
            w84=> c1_n4_w84, 
            w85=> c1_n4_w85, 
            w86=> c1_n4_w86, 
            w87=> c1_n4_w87, 
            w88=> c1_n4_w88, 
            w89=> c1_n4_w89, 
            w90=> c1_n4_w90, 
            w91=> c1_n4_w91, 
            w92=> c1_n4_w92, 
            w93=> c1_n4_w93, 
            w94=> c1_n4_w94, 
            w95=> c1_n4_w95, 
            w96=> c1_n4_w96, 
            w97=> c1_n4_w97, 
            w98=> c1_n4_w98, 
            w99=> c1_n4_w99, 
            w100=> c1_n4_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n5_w1, 
            w2=> c1_n5_w2, 
            w3=> c1_n5_w3, 
            w4=> c1_n5_w4, 
            w5=> c1_n5_w5, 
            w6=> c1_n5_w6, 
            w7=> c1_n5_w7, 
            w8=> c1_n5_w8, 
            w9=> c1_n5_w9, 
            w10=> c1_n5_w10, 
            w11=> c1_n5_w11, 
            w12=> c1_n5_w12, 
            w13=> c1_n5_w13, 
            w14=> c1_n5_w14, 
            w15=> c1_n5_w15, 
            w16=> c1_n5_w16, 
            w17=> c1_n5_w17, 
            w18=> c1_n5_w18, 
            w19=> c1_n5_w19, 
            w20=> c1_n5_w20, 
            w21=> c1_n5_w21, 
            w22=> c1_n5_w22, 
            w23=> c1_n5_w23, 
            w24=> c1_n5_w24, 
            w25=> c1_n5_w25, 
            w26=> c1_n5_w26, 
            w27=> c1_n5_w27, 
            w28=> c1_n5_w28, 
            w29=> c1_n5_w29, 
            w30=> c1_n5_w30, 
            w31=> c1_n5_w31, 
            w32=> c1_n5_w32, 
            w33=> c1_n5_w33, 
            w34=> c1_n5_w34, 
            w35=> c1_n5_w35, 
            w36=> c1_n5_w36, 
            w37=> c1_n5_w37, 
            w38=> c1_n5_w38, 
            w39=> c1_n5_w39, 
            w40=> c1_n5_w40, 
            w41=> c1_n5_w41, 
            w42=> c1_n5_w42, 
            w43=> c1_n5_w43, 
            w44=> c1_n5_w44, 
            w45=> c1_n5_w45, 
            w46=> c1_n5_w46, 
            w47=> c1_n5_w47, 
            w48=> c1_n5_w48, 
            w49=> c1_n5_w49, 
            w50=> c1_n5_w50, 
            w51=> c1_n5_w51, 
            w52=> c1_n5_w52, 
            w53=> c1_n5_w53, 
            w54=> c1_n5_w54, 
            w55=> c1_n5_w55, 
            w56=> c1_n5_w56, 
            w57=> c1_n5_w57, 
            w58=> c1_n5_w58, 
            w59=> c1_n5_w59, 
            w60=> c1_n5_w60, 
            w61=> c1_n5_w61, 
            w62=> c1_n5_w62, 
            w63=> c1_n5_w63, 
            w64=> c1_n5_w64, 
            w65=> c1_n5_w65, 
            w66=> c1_n5_w66, 
            w67=> c1_n5_w67, 
            w68=> c1_n5_w68, 
            w69=> c1_n5_w69, 
            w70=> c1_n5_w70, 
            w71=> c1_n5_w71, 
            w72=> c1_n5_w72, 
            w73=> c1_n5_w73, 
            w74=> c1_n5_w74, 
            w75=> c1_n5_w75, 
            w76=> c1_n5_w76, 
            w77=> c1_n5_w77, 
            w78=> c1_n5_w78, 
            w79=> c1_n5_w79, 
            w80=> c1_n5_w80, 
            w81=> c1_n5_w81, 
            w82=> c1_n5_w82, 
            w83=> c1_n5_w83, 
            w84=> c1_n5_w84, 
            w85=> c1_n5_w85, 
            w86=> c1_n5_w86, 
            w87=> c1_n5_w87, 
            w88=> c1_n5_w88, 
            w89=> c1_n5_w89, 
            w90=> c1_n5_w90, 
            w91=> c1_n5_w91, 
            w92=> c1_n5_w92, 
            w93=> c1_n5_w93, 
            w94=> c1_n5_w94, 
            w95=> c1_n5_w95, 
            w96=> c1_n5_w96, 
            w97=> c1_n5_w97, 
            w98=> c1_n5_w98, 
            w99=> c1_n5_w99, 
            w100=> c1_n5_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n6_w1, 
            w2=> c1_n6_w2, 
            w3=> c1_n6_w3, 
            w4=> c1_n6_w4, 
            w5=> c1_n6_w5, 
            w6=> c1_n6_w6, 
            w7=> c1_n6_w7, 
            w8=> c1_n6_w8, 
            w9=> c1_n6_w9, 
            w10=> c1_n6_w10, 
            w11=> c1_n6_w11, 
            w12=> c1_n6_w12, 
            w13=> c1_n6_w13, 
            w14=> c1_n6_w14, 
            w15=> c1_n6_w15, 
            w16=> c1_n6_w16, 
            w17=> c1_n6_w17, 
            w18=> c1_n6_w18, 
            w19=> c1_n6_w19, 
            w20=> c1_n6_w20, 
            w21=> c1_n6_w21, 
            w22=> c1_n6_w22, 
            w23=> c1_n6_w23, 
            w24=> c1_n6_w24, 
            w25=> c1_n6_w25, 
            w26=> c1_n6_w26, 
            w27=> c1_n6_w27, 
            w28=> c1_n6_w28, 
            w29=> c1_n6_w29, 
            w30=> c1_n6_w30, 
            w31=> c1_n6_w31, 
            w32=> c1_n6_w32, 
            w33=> c1_n6_w33, 
            w34=> c1_n6_w34, 
            w35=> c1_n6_w35, 
            w36=> c1_n6_w36, 
            w37=> c1_n6_w37, 
            w38=> c1_n6_w38, 
            w39=> c1_n6_w39, 
            w40=> c1_n6_w40, 
            w41=> c1_n6_w41, 
            w42=> c1_n6_w42, 
            w43=> c1_n6_w43, 
            w44=> c1_n6_w44, 
            w45=> c1_n6_w45, 
            w46=> c1_n6_w46, 
            w47=> c1_n6_w47, 
            w48=> c1_n6_w48, 
            w49=> c1_n6_w49, 
            w50=> c1_n6_w50, 
            w51=> c1_n6_w51, 
            w52=> c1_n6_w52, 
            w53=> c1_n6_w53, 
            w54=> c1_n6_w54, 
            w55=> c1_n6_w55, 
            w56=> c1_n6_w56, 
            w57=> c1_n6_w57, 
            w58=> c1_n6_w58, 
            w59=> c1_n6_w59, 
            w60=> c1_n6_w60, 
            w61=> c1_n6_w61, 
            w62=> c1_n6_w62, 
            w63=> c1_n6_w63, 
            w64=> c1_n6_w64, 
            w65=> c1_n6_w65, 
            w66=> c1_n6_w66, 
            w67=> c1_n6_w67, 
            w68=> c1_n6_w68, 
            w69=> c1_n6_w69, 
            w70=> c1_n6_w70, 
            w71=> c1_n6_w71, 
            w72=> c1_n6_w72, 
            w73=> c1_n6_w73, 
            w74=> c1_n6_w74, 
            w75=> c1_n6_w75, 
            w76=> c1_n6_w76, 
            w77=> c1_n6_w77, 
            w78=> c1_n6_w78, 
            w79=> c1_n6_w79, 
            w80=> c1_n6_w80, 
            w81=> c1_n6_w81, 
            w82=> c1_n6_w82, 
            w83=> c1_n6_w83, 
            w84=> c1_n6_w84, 
            w85=> c1_n6_w85, 
            w86=> c1_n6_w86, 
            w87=> c1_n6_w87, 
            w88=> c1_n6_w88, 
            w89=> c1_n6_w89, 
            w90=> c1_n6_w90, 
            w91=> c1_n6_w91, 
            w92=> c1_n6_w92, 
            w93=> c1_n6_w93, 
            w94=> c1_n6_w94, 
            w95=> c1_n6_w95, 
            w96=> c1_n6_w96, 
            w97=> c1_n6_w97, 
            w98=> c1_n6_w98, 
            w99=> c1_n6_w99, 
            w100=> c1_n6_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n7_w1, 
            w2=> c1_n7_w2, 
            w3=> c1_n7_w3, 
            w4=> c1_n7_w4, 
            w5=> c1_n7_w5, 
            w6=> c1_n7_w6, 
            w7=> c1_n7_w7, 
            w8=> c1_n7_w8, 
            w9=> c1_n7_w9, 
            w10=> c1_n7_w10, 
            w11=> c1_n7_w11, 
            w12=> c1_n7_w12, 
            w13=> c1_n7_w13, 
            w14=> c1_n7_w14, 
            w15=> c1_n7_w15, 
            w16=> c1_n7_w16, 
            w17=> c1_n7_w17, 
            w18=> c1_n7_w18, 
            w19=> c1_n7_w19, 
            w20=> c1_n7_w20, 
            w21=> c1_n7_w21, 
            w22=> c1_n7_w22, 
            w23=> c1_n7_w23, 
            w24=> c1_n7_w24, 
            w25=> c1_n7_w25, 
            w26=> c1_n7_w26, 
            w27=> c1_n7_w27, 
            w28=> c1_n7_w28, 
            w29=> c1_n7_w29, 
            w30=> c1_n7_w30, 
            w31=> c1_n7_w31, 
            w32=> c1_n7_w32, 
            w33=> c1_n7_w33, 
            w34=> c1_n7_w34, 
            w35=> c1_n7_w35, 
            w36=> c1_n7_w36, 
            w37=> c1_n7_w37, 
            w38=> c1_n7_w38, 
            w39=> c1_n7_w39, 
            w40=> c1_n7_w40, 
            w41=> c1_n7_w41, 
            w42=> c1_n7_w42, 
            w43=> c1_n7_w43, 
            w44=> c1_n7_w44, 
            w45=> c1_n7_w45, 
            w46=> c1_n7_w46, 
            w47=> c1_n7_w47, 
            w48=> c1_n7_w48, 
            w49=> c1_n7_w49, 
            w50=> c1_n7_w50, 
            w51=> c1_n7_w51, 
            w52=> c1_n7_w52, 
            w53=> c1_n7_w53, 
            w54=> c1_n7_w54, 
            w55=> c1_n7_w55, 
            w56=> c1_n7_w56, 
            w57=> c1_n7_w57, 
            w58=> c1_n7_w58, 
            w59=> c1_n7_w59, 
            w60=> c1_n7_w60, 
            w61=> c1_n7_w61, 
            w62=> c1_n7_w62, 
            w63=> c1_n7_w63, 
            w64=> c1_n7_w64, 
            w65=> c1_n7_w65, 
            w66=> c1_n7_w66, 
            w67=> c1_n7_w67, 
            w68=> c1_n7_w68, 
            w69=> c1_n7_w69, 
            w70=> c1_n7_w70, 
            w71=> c1_n7_w71, 
            w72=> c1_n7_w72, 
            w73=> c1_n7_w73, 
            w74=> c1_n7_w74, 
            w75=> c1_n7_w75, 
            w76=> c1_n7_w76, 
            w77=> c1_n7_w77, 
            w78=> c1_n7_w78, 
            w79=> c1_n7_w79, 
            w80=> c1_n7_w80, 
            w81=> c1_n7_w81, 
            w82=> c1_n7_w82, 
            w83=> c1_n7_w83, 
            w84=> c1_n7_w84, 
            w85=> c1_n7_w85, 
            w86=> c1_n7_w86, 
            w87=> c1_n7_w87, 
            w88=> c1_n7_w88, 
            w89=> c1_n7_w89, 
            w90=> c1_n7_w90, 
            w91=> c1_n7_w91, 
            w92=> c1_n7_w92, 
            w93=> c1_n7_w93, 
            w94=> c1_n7_w94, 
            w95=> c1_n7_w95, 
            w96=> c1_n7_w96, 
            w97=> c1_n7_w97, 
            w98=> c1_n7_w98, 
            w99=> c1_n7_w99, 
            w100=> c1_n7_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n8_w1, 
            w2=> c1_n8_w2, 
            w3=> c1_n8_w3, 
            w4=> c1_n8_w4, 
            w5=> c1_n8_w5, 
            w6=> c1_n8_w6, 
            w7=> c1_n8_w7, 
            w8=> c1_n8_w8, 
            w9=> c1_n8_w9, 
            w10=> c1_n8_w10, 
            w11=> c1_n8_w11, 
            w12=> c1_n8_w12, 
            w13=> c1_n8_w13, 
            w14=> c1_n8_w14, 
            w15=> c1_n8_w15, 
            w16=> c1_n8_w16, 
            w17=> c1_n8_w17, 
            w18=> c1_n8_w18, 
            w19=> c1_n8_w19, 
            w20=> c1_n8_w20, 
            w21=> c1_n8_w21, 
            w22=> c1_n8_w22, 
            w23=> c1_n8_w23, 
            w24=> c1_n8_w24, 
            w25=> c1_n8_w25, 
            w26=> c1_n8_w26, 
            w27=> c1_n8_w27, 
            w28=> c1_n8_w28, 
            w29=> c1_n8_w29, 
            w30=> c1_n8_w30, 
            w31=> c1_n8_w31, 
            w32=> c1_n8_w32, 
            w33=> c1_n8_w33, 
            w34=> c1_n8_w34, 
            w35=> c1_n8_w35, 
            w36=> c1_n8_w36, 
            w37=> c1_n8_w37, 
            w38=> c1_n8_w38, 
            w39=> c1_n8_w39, 
            w40=> c1_n8_w40, 
            w41=> c1_n8_w41, 
            w42=> c1_n8_w42, 
            w43=> c1_n8_w43, 
            w44=> c1_n8_w44, 
            w45=> c1_n8_w45, 
            w46=> c1_n8_w46, 
            w47=> c1_n8_w47, 
            w48=> c1_n8_w48, 
            w49=> c1_n8_w49, 
            w50=> c1_n8_w50, 
            w51=> c1_n8_w51, 
            w52=> c1_n8_w52, 
            w53=> c1_n8_w53, 
            w54=> c1_n8_w54, 
            w55=> c1_n8_w55, 
            w56=> c1_n8_w56, 
            w57=> c1_n8_w57, 
            w58=> c1_n8_w58, 
            w59=> c1_n8_w59, 
            w60=> c1_n8_w60, 
            w61=> c1_n8_w61, 
            w62=> c1_n8_w62, 
            w63=> c1_n8_w63, 
            w64=> c1_n8_w64, 
            w65=> c1_n8_w65, 
            w66=> c1_n8_w66, 
            w67=> c1_n8_w67, 
            w68=> c1_n8_w68, 
            w69=> c1_n8_w69, 
            w70=> c1_n8_w70, 
            w71=> c1_n8_w71, 
            w72=> c1_n8_w72, 
            w73=> c1_n8_w73, 
            w74=> c1_n8_w74, 
            w75=> c1_n8_w75, 
            w76=> c1_n8_w76, 
            w77=> c1_n8_w77, 
            w78=> c1_n8_w78, 
            w79=> c1_n8_w79, 
            w80=> c1_n8_w80, 
            w81=> c1_n8_w81, 
            w82=> c1_n8_w82, 
            w83=> c1_n8_w83, 
            w84=> c1_n8_w84, 
            w85=> c1_n8_w85, 
            w86=> c1_n8_w86, 
            w87=> c1_n8_w87, 
            w88=> c1_n8_w88, 
            w89=> c1_n8_w89, 
            w90=> c1_n8_w90, 
            w91=> c1_n8_w91, 
            w92=> c1_n8_w92, 
            w93=> c1_n8_w93, 
            w94=> c1_n8_w94, 
            w95=> c1_n8_w95, 
            w96=> c1_n8_w96, 
            w97=> c1_n8_w97, 
            w98=> c1_n8_w98, 
            w99=> c1_n8_w99, 
            w100=> c1_n8_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n9_w1, 
            w2=> c1_n9_w2, 
            w3=> c1_n9_w3, 
            w4=> c1_n9_w4, 
            w5=> c1_n9_w5, 
            w6=> c1_n9_w6, 
            w7=> c1_n9_w7, 
            w8=> c1_n9_w8, 
            w9=> c1_n9_w9, 
            w10=> c1_n9_w10, 
            w11=> c1_n9_w11, 
            w12=> c1_n9_w12, 
            w13=> c1_n9_w13, 
            w14=> c1_n9_w14, 
            w15=> c1_n9_w15, 
            w16=> c1_n9_w16, 
            w17=> c1_n9_w17, 
            w18=> c1_n9_w18, 
            w19=> c1_n9_w19, 
            w20=> c1_n9_w20, 
            w21=> c1_n9_w21, 
            w22=> c1_n9_w22, 
            w23=> c1_n9_w23, 
            w24=> c1_n9_w24, 
            w25=> c1_n9_w25, 
            w26=> c1_n9_w26, 
            w27=> c1_n9_w27, 
            w28=> c1_n9_w28, 
            w29=> c1_n9_w29, 
            w30=> c1_n9_w30, 
            w31=> c1_n9_w31, 
            w32=> c1_n9_w32, 
            w33=> c1_n9_w33, 
            w34=> c1_n9_w34, 
            w35=> c1_n9_w35, 
            w36=> c1_n9_w36, 
            w37=> c1_n9_w37, 
            w38=> c1_n9_w38, 
            w39=> c1_n9_w39, 
            w40=> c1_n9_w40, 
            w41=> c1_n9_w41, 
            w42=> c1_n9_w42, 
            w43=> c1_n9_w43, 
            w44=> c1_n9_w44, 
            w45=> c1_n9_w45, 
            w46=> c1_n9_w46, 
            w47=> c1_n9_w47, 
            w48=> c1_n9_w48, 
            w49=> c1_n9_w49, 
            w50=> c1_n9_w50, 
            w51=> c1_n9_w51, 
            w52=> c1_n9_w52, 
            w53=> c1_n9_w53, 
            w54=> c1_n9_w54, 
            w55=> c1_n9_w55, 
            w56=> c1_n9_w56, 
            w57=> c1_n9_w57, 
            w58=> c1_n9_w58, 
            w59=> c1_n9_w59, 
            w60=> c1_n9_w60, 
            w61=> c1_n9_w61, 
            w62=> c1_n9_w62, 
            w63=> c1_n9_w63, 
            w64=> c1_n9_w64, 
            w65=> c1_n9_w65, 
            w66=> c1_n9_w66, 
            w67=> c1_n9_w67, 
            w68=> c1_n9_w68, 
            w69=> c1_n9_w69, 
            w70=> c1_n9_w70, 
            w71=> c1_n9_w71, 
            w72=> c1_n9_w72, 
            w73=> c1_n9_w73, 
            w74=> c1_n9_w74, 
            w75=> c1_n9_w75, 
            w76=> c1_n9_w76, 
            w77=> c1_n9_w77, 
            w78=> c1_n9_w78, 
            w79=> c1_n9_w79, 
            w80=> c1_n9_w80, 
            w81=> c1_n9_w81, 
            w82=> c1_n9_w82, 
            w83=> c1_n9_w83, 
            w84=> c1_n9_w84, 
            w85=> c1_n9_w85, 
            w86=> c1_n9_w86, 
            w87=> c1_n9_w87, 
            w88=> c1_n9_w88, 
            w89=> c1_n9_w89, 
            w90=> c1_n9_w90, 
            w91=> c1_n9_w91, 
            w92=> c1_n9_w92, 
            w93=> c1_n9_w93, 
            w94=> c1_n9_w94, 
            w95=> c1_n9_w95, 
            w96=> c1_n9_w96, 
            w97=> c1_n9_w97, 
            w98=> c1_n9_w98, 
            w99=> c1_n9_w99, 
            w100=> c1_n9_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n9_y
   );           
            
neuron_inst_10: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n10_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n10_w1, 
            w2=> c1_n10_w2, 
            w3=> c1_n10_w3, 
            w4=> c1_n10_w4, 
            w5=> c1_n10_w5, 
            w6=> c1_n10_w6, 
            w7=> c1_n10_w7, 
            w8=> c1_n10_w8, 
            w9=> c1_n10_w9, 
            w10=> c1_n10_w10, 
            w11=> c1_n10_w11, 
            w12=> c1_n10_w12, 
            w13=> c1_n10_w13, 
            w14=> c1_n10_w14, 
            w15=> c1_n10_w15, 
            w16=> c1_n10_w16, 
            w17=> c1_n10_w17, 
            w18=> c1_n10_w18, 
            w19=> c1_n10_w19, 
            w20=> c1_n10_w20, 
            w21=> c1_n10_w21, 
            w22=> c1_n10_w22, 
            w23=> c1_n10_w23, 
            w24=> c1_n10_w24, 
            w25=> c1_n10_w25, 
            w26=> c1_n10_w26, 
            w27=> c1_n10_w27, 
            w28=> c1_n10_w28, 
            w29=> c1_n10_w29, 
            w30=> c1_n10_w30, 
            w31=> c1_n10_w31, 
            w32=> c1_n10_w32, 
            w33=> c1_n10_w33, 
            w34=> c1_n10_w34, 
            w35=> c1_n10_w35, 
            w36=> c1_n10_w36, 
            w37=> c1_n10_w37, 
            w38=> c1_n10_w38, 
            w39=> c1_n10_w39, 
            w40=> c1_n10_w40, 
            w41=> c1_n10_w41, 
            w42=> c1_n10_w42, 
            w43=> c1_n10_w43, 
            w44=> c1_n10_w44, 
            w45=> c1_n10_w45, 
            w46=> c1_n10_w46, 
            w47=> c1_n10_w47, 
            w48=> c1_n10_w48, 
            w49=> c1_n10_w49, 
            w50=> c1_n10_w50, 
            w51=> c1_n10_w51, 
            w52=> c1_n10_w52, 
            w53=> c1_n10_w53, 
            w54=> c1_n10_w54, 
            w55=> c1_n10_w55, 
            w56=> c1_n10_w56, 
            w57=> c1_n10_w57, 
            w58=> c1_n10_w58, 
            w59=> c1_n10_w59, 
            w60=> c1_n10_w60, 
            w61=> c1_n10_w61, 
            w62=> c1_n10_w62, 
            w63=> c1_n10_w63, 
            w64=> c1_n10_w64, 
            w65=> c1_n10_w65, 
            w66=> c1_n10_w66, 
            w67=> c1_n10_w67, 
            w68=> c1_n10_w68, 
            w69=> c1_n10_w69, 
            w70=> c1_n10_w70, 
            w71=> c1_n10_w71, 
            w72=> c1_n10_w72, 
            w73=> c1_n10_w73, 
            w74=> c1_n10_w74, 
            w75=> c1_n10_w75, 
            w76=> c1_n10_w76, 
            w77=> c1_n10_w77, 
            w78=> c1_n10_w78, 
            w79=> c1_n10_w79, 
            w80=> c1_n10_w80, 
            w81=> c1_n10_w81, 
            w82=> c1_n10_w82, 
            w83=> c1_n10_w83, 
            w84=> c1_n10_w84, 
            w85=> c1_n10_w85, 
            w86=> c1_n10_w86, 
            w87=> c1_n10_w87, 
            w88=> c1_n10_w88, 
            w89=> c1_n10_w89, 
            w90=> c1_n10_w90, 
            w91=> c1_n10_w91, 
            w92=> c1_n10_w92, 
            w93=> c1_n10_w93, 
            w94=> c1_n10_w94, 
            w95=> c1_n10_w95, 
            w96=> c1_n10_w96, 
            w97=> c1_n10_w97, 
            w98=> c1_n10_w98, 
            w99=> c1_n10_w99, 
            w100=> c1_n10_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n10_y
   );           
            
neuron_inst_11: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n11_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n11_w1, 
            w2=> c1_n11_w2, 
            w3=> c1_n11_w3, 
            w4=> c1_n11_w4, 
            w5=> c1_n11_w5, 
            w6=> c1_n11_w6, 
            w7=> c1_n11_w7, 
            w8=> c1_n11_w8, 
            w9=> c1_n11_w9, 
            w10=> c1_n11_w10, 
            w11=> c1_n11_w11, 
            w12=> c1_n11_w12, 
            w13=> c1_n11_w13, 
            w14=> c1_n11_w14, 
            w15=> c1_n11_w15, 
            w16=> c1_n11_w16, 
            w17=> c1_n11_w17, 
            w18=> c1_n11_w18, 
            w19=> c1_n11_w19, 
            w20=> c1_n11_w20, 
            w21=> c1_n11_w21, 
            w22=> c1_n11_w22, 
            w23=> c1_n11_w23, 
            w24=> c1_n11_w24, 
            w25=> c1_n11_w25, 
            w26=> c1_n11_w26, 
            w27=> c1_n11_w27, 
            w28=> c1_n11_w28, 
            w29=> c1_n11_w29, 
            w30=> c1_n11_w30, 
            w31=> c1_n11_w31, 
            w32=> c1_n11_w32, 
            w33=> c1_n11_w33, 
            w34=> c1_n11_w34, 
            w35=> c1_n11_w35, 
            w36=> c1_n11_w36, 
            w37=> c1_n11_w37, 
            w38=> c1_n11_w38, 
            w39=> c1_n11_w39, 
            w40=> c1_n11_w40, 
            w41=> c1_n11_w41, 
            w42=> c1_n11_w42, 
            w43=> c1_n11_w43, 
            w44=> c1_n11_w44, 
            w45=> c1_n11_w45, 
            w46=> c1_n11_w46, 
            w47=> c1_n11_w47, 
            w48=> c1_n11_w48, 
            w49=> c1_n11_w49, 
            w50=> c1_n11_w50, 
            w51=> c1_n11_w51, 
            w52=> c1_n11_w52, 
            w53=> c1_n11_w53, 
            w54=> c1_n11_w54, 
            w55=> c1_n11_w55, 
            w56=> c1_n11_w56, 
            w57=> c1_n11_w57, 
            w58=> c1_n11_w58, 
            w59=> c1_n11_w59, 
            w60=> c1_n11_w60, 
            w61=> c1_n11_w61, 
            w62=> c1_n11_w62, 
            w63=> c1_n11_w63, 
            w64=> c1_n11_w64, 
            w65=> c1_n11_w65, 
            w66=> c1_n11_w66, 
            w67=> c1_n11_w67, 
            w68=> c1_n11_w68, 
            w69=> c1_n11_w69, 
            w70=> c1_n11_w70, 
            w71=> c1_n11_w71, 
            w72=> c1_n11_w72, 
            w73=> c1_n11_w73, 
            w74=> c1_n11_w74, 
            w75=> c1_n11_w75, 
            w76=> c1_n11_w76, 
            w77=> c1_n11_w77, 
            w78=> c1_n11_w78, 
            w79=> c1_n11_w79, 
            w80=> c1_n11_w80, 
            w81=> c1_n11_w81, 
            w82=> c1_n11_w82, 
            w83=> c1_n11_w83, 
            w84=> c1_n11_w84, 
            w85=> c1_n11_w85, 
            w86=> c1_n11_w86, 
            w87=> c1_n11_w87, 
            w88=> c1_n11_w88, 
            w89=> c1_n11_w89, 
            w90=> c1_n11_w90, 
            w91=> c1_n11_w91, 
            w92=> c1_n11_w92, 
            w93=> c1_n11_w93, 
            w94=> c1_n11_w94, 
            w95=> c1_n11_w95, 
            w96=> c1_n11_w96, 
            w97=> c1_n11_w97, 
            w98=> c1_n11_w98, 
            w99=> c1_n11_w99, 
            w100=> c1_n11_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n11_y
   );           
            
neuron_inst_12: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n12_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n12_w1, 
            w2=> c1_n12_w2, 
            w3=> c1_n12_w3, 
            w4=> c1_n12_w4, 
            w5=> c1_n12_w5, 
            w6=> c1_n12_w6, 
            w7=> c1_n12_w7, 
            w8=> c1_n12_w8, 
            w9=> c1_n12_w9, 
            w10=> c1_n12_w10, 
            w11=> c1_n12_w11, 
            w12=> c1_n12_w12, 
            w13=> c1_n12_w13, 
            w14=> c1_n12_w14, 
            w15=> c1_n12_w15, 
            w16=> c1_n12_w16, 
            w17=> c1_n12_w17, 
            w18=> c1_n12_w18, 
            w19=> c1_n12_w19, 
            w20=> c1_n12_w20, 
            w21=> c1_n12_w21, 
            w22=> c1_n12_w22, 
            w23=> c1_n12_w23, 
            w24=> c1_n12_w24, 
            w25=> c1_n12_w25, 
            w26=> c1_n12_w26, 
            w27=> c1_n12_w27, 
            w28=> c1_n12_w28, 
            w29=> c1_n12_w29, 
            w30=> c1_n12_w30, 
            w31=> c1_n12_w31, 
            w32=> c1_n12_w32, 
            w33=> c1_n12_w33, 
            w34=> c1_n12_w34, 
            w35=> c1_n12_w35, 
            w36=> c1_n12_w36, 
            w37=> c1_n12_w37, 
            w38=> c1_n12_w38, 
            w39=> c1_n12_w39, 
            w40=> c1_n12_w40, 
            w41=> c1_n12_w41, 
            w42=> c1_n12_w42, 
            w43=> c1_n12_w43, 
            w44=> c1_n12_w44, 
            w45=> c1_n12_w45, 
            w46=> c1_n12_w46, 
            w47=> c1_n12_w47, 
            w48=> c1_n12_w48, 
            w49=> c1_n12_w49, 
            w50=> c1_n12_w50, 
            w51=> c1_n12_w51, 
            w52=> c1_n12_w52, 
            w53=> c1_n12_w53, 
            w54=> c1_n12_w54, 
            w55=> c1_n12_w55, 
            w56=> c1_n12_w56, 
            w57=> c1_n12_w57, 
            w58=> c1_n12_w58, 
            w59=> c1_n12_w59, 
            w60=> c1_n12_w60, 
            w61=> c1_n12_w61, 
            w62=> c1_n12_w62, 
            w63=> c1_n12_w63, 
            w64=> c1_n12_w64, 
            w65=> c1_n12_w65, 
            w66=> c1_n12_w66, 
            w67=> c1_n12_w67, 
            w68=> c1_n12_w68, 
            w69=> c1_n12_w69, 
            w70=> c1_n12_w70, 
            w71=> c1_n12_w71, 
            w72=> c1_n12_w72, 
            w73=> c1_n12_w73, 
            w74=> c1_n12_w74, 
            w75=> c1_n12_w75, 
            w76=> c1_n12_w76, 
            w77=> c1_n12_w77, 
            w78=> c1_n12_w78, 
            w79=> c1_n12_w79, 
            w80=> c1_n12_w80, 
            w81=> c1_n12_w81, 
            w82=> c1_n12_w82, 
            w83=> c1_n12_w83, 
            w84=> c1_n12_w84, 
            w85=> c1_n12_w85, 
            w86=> c1_n12_w86, 
            w87=> c1_n12_w87, 
            w88=> c1_n12_w88, 
            w89=> c1_n12_w89, 
            w90=> c1_n12_w90, 
            w91=> c1_n12_w91, 
            w92=> c1_n12_w92, 
            w93=> c1_n12_w93, 
            w94=> c1_n12_w94, 
            w95=> c1_n12_w95, 
            w96=> c1_n12_w96, 
            w97=> c1_n12_w97, 
            w98=> c1_n12_w98, 
            w99=> c1_n12_w99, 
            w100=> c1_n12_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n12_y
   );           
            
neuron_inst_13: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n13_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n13_w1, 
            w2=> c1_n13_w2, 
            w3=> c1_n13_w3, 
            w4=> c1_n13_w4, 
            w5=> c1_n13_w5, 
            w6=> c1_n13_w6, 
            w7=> c1_n13_w7, 
            w8=> c1_n13_w8, 
            w9=> c1_n13_w9, 
            w10=> c1_n13_w10, 
            w11=> c1_n13_w11, 
            w12=> c1_n13_w12, 
            w13=> c1_n13_w13, 
            w14=> c1_n13_w14, 
            w15=> c1_n13_w15, 
            w16=> c1_n13_w16, 
            w17=> c1_n13_w17, 
            w18=> c1_n13_w18, 
            w19=> c1_n13_w19, 
            w20=> c1_n13_w20, 
            w21=> c1_n13_w21, 
            w22=> c1_n13_w22, 
            w23=> c1_n13_w23, 
            w24=> c1_n13_w24, 
            w25=> c1_n13_w25, 
            w26=> c1_n13_w26, 
            w27=> c1_n13_w27, 
            w28=> c1_n13_w28, 
            w29=> c1_n13_w29, 
            w30=> c1_n13_w30, 
            w31=> c1_n13_w31, 
            w32=> c1_n13_w32, 
            w33=> c1_n13_w33, 
            w34=> c1_n13_w34, 
            w35=> c1_n13_w35, 
            w36=> c1_n13_w36, 
            w37=> c1_n13_w37, 
            w38=> c1_n13_w38, 
            w39=> c1_n13_w39, 
            w40=> c1_n13_w40, 
            w41=> c1_n13_w41, 
            w42=> c1_n13_w42, 
            w43=> c1_n13_w43, 
            w44=> c1_n13_w44, 
            w45=> c1_n13_w45, 
            w46=> c1_n13_w46, 
            w47=> c1_n13_w47, 
            w48=> c1_n13_w48, 
            w49=> c1_n13_w49, 
            w50=> c1_n13_w50, 
            w51=> c1_n13_w51, 
            w52=> c1_n13_w52, 
            w53=> c1_n13_w53, 
            w54=> c1_n13_w54, 
            w55=> c1_n13_w55, 
            w56=> c1_n13_w56, 
            w57=> c1_n13_w57, 
            w58=> c1_n13_w58, 
            w59=> c1_n13_w59, 
            w60=> c1_n13_w60, 
            w61=> c1_n13_w61, 
            w62=> c1_n13_w62, 
            w63=> c1_n13_w63, 
            w64=> c1_n13_w64, 
            w65=> c1_n13_w65, 
            w66=> c1_n13_w66, 
            w67=> c1_n13_w67, 
            w68=> c1_n13_w68, 
            w69=> c1_n13_w69, 
            w70=> c1_n13_w70, 
            w71=> c1_n13_w71, 
            w72=> c1_n13_w72, 
            w73=> c1_n13_w73, 
            w74=> c1_n13_w74, 
            w75=> c1_n13_w75, 
            w76=> c1_n13_w76, 
            w77=> c1_n13_w77, 
            w78=> c1_n13_w78, 
            w79=> c1_n13_w79, 
            w80=> c1_n13_w80, 
            w81=> c1_n13_w81, 
            w82=> c1_n13_w82, 
            w83=> c1_n13_w83, 
            w84=> c1_n13_w84, 
            w85=> c1_n13_w85, 
            w86=> c1_n13_w86, 
            w87=> c1_n13_w87, 
            w88=> c1_n13_w88, 
            w89=> c1_n13_w89, 
            w90=> c1_n13_w90, 
            w91=> c1_n13_w91, 
            w92=> c1_n13_w92, 
            w93=> c1_n13_w93, 
            w94=> c1_n13_w94, 
            w95=> c1_n13_w95, 
            w96=> c1_n13_w96, 
            w97=> c1_n13_w97, 
            w98=> c1_n13_w98, 
            w99=> c1_n13_w99, 
            w100=> c1_n13_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n13_y
   );           
            
neuron_inst_14: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n14_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n14_w1, 
            w2=> c1_n14_w2, 
            w3=> c1_n14_w3, 
            w4=> c1_n14_w4, 
            w5=> c1_n14_w5, 
            w6=> c1_n14_w6, 
            w7=> c1_n14_w7, 
            w8=> c1_n14_w8, 
            w9=> c1_n14_w9, 
            w10=> c1_n14_w10, 
            w11=> c1_n14_w11, 
            w12=> c1_n14_w12, 
            w13=> c1_n14_w13, 
            w14=> c1_n14_w14, 
            w15=> c1_n14_w15, 
            w16=> c1_n14_w16, 
            w17=> c1_n14_w17, 
            w18=> c1_n14_w18, 
            w19=> c1_n14_w19, 
            w20=> c1_n14_w20, 
            w21=> c1_n14_w21, 
            w22=> c1_n14_w22, 
            w23=> c1_n14_w23, 
            w24=> c1_n14_w24, 
            w25=> c1_n14_w25, 
            w26=> c1_n14_w26, 
            w27=> c1_n14_w27, 
            w28=> c1_n14_w28, 
            w29=> c1_n14_w29, 
            w30=> c1_n14_w30, 
            w31=> c1_n14_w31, 
            w32=> c1_n14_w32, 
            w33=> c1_n14_w33, 
            w34=> c1_n14_w34, 
            w35=> c1_n14_w35, 
            w36=> c1_n14_w36, 
            w37=> c1_n14_w37, 
            w38=> c1_n14_w38, 
            w39=> c1_n14_w39, 
            w40=> c1_n14_w40, 
            w41=> c1_n14_w41, 
            w42=> c1_n14_w42, 
            w43=> c1_n14_w43, 
            w44=> c1_n14_w44, 
            w45=> c1_n14_w45, 
            w46=> c1_n14_w46, 
            w47=> c1_n14_w47, 
            w48=> c1_n14_w48, 
            w49=> c1_n14_w49, 
            w50=> c1_n14_w50, 
            w51=> c1_n14_w51, 
            w52=> c1_n14_w52, 
            w53=> c1_n14_w53, 
            w54=> c1_n14_w54, 
            w55=> c1_n14_w55, 
            w56=> c1_n14_w56, 
            w57=> c1_n14_w57, 
            w58=> c1_n14_w58, 
            w59=> c1_n14_w59, 
            w60=> c1_n14_w60, 
            w61=> c1_n14_w61, 
            w62=> c1_n14_w62, 
            w63=> c1_n14_w63, 
            w64=> c1_n14_w64, 
            w65=> c1_n14_w65, 
            w66=> c1_n14_w66, 
            w67=> c1_n14_w67, 
            w68=> c1_n14_w68, 
            w69=> c1_n14_w69, 
            w70=> c1_n14_w70, 
            w71=> c1_n14_w71, 
            w72=> c1_n14_w72, 
            w73=> c1_n14_w73, 
            w74=> c1_n14_w74, 
            w75=> c1_n14_w75, 
            w76=> c1_n14_w76, 
            w77=> c1_n14_w77, 
            w78=> c1_n14_w78, 
            w79=> c1_n14_w79, 
            w80=> c1_n14_w80, 
            w81=> c1_n14_w81, 
            w82=> c1_n14_w82, 
            w83=> c1_n14_w83, 
            w84=> c1_n14_w84, 
            w85=> c1_n14_w85, 
            w86=> c1_n14_w86, 
            w87=> c1_n14_w87, 
            w88=> c1_n14_w88, 
            w89=> c1_n14_w89, 
            w90=> c1_n14_w90, 
            w91=> c1_n14_w91, 
            w92=> c1_n14_w92, 
            w93=> c1_n14_w93, 
            w94=> c1_n14_w94, 
            w95=> c1_n14_w95, 
            w96=> c1_n14_w96, 
            w97=> c1_n14_w97, 
            w98=> c1_n14_w98, 
            w99=> c1_n14_w99, 
            w100=> c1_n14_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n14_y
   );           
            
neuron_inst_15: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n15_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n15_w1, 
            w2=> c1_n15_w2, 
            w3=> c1_n15_w3, 
            w4=> c1_n15_w4, 
            w5=> c1_n15_w5, 
            w6=> c1_n15_w6, 
            w7=> c1_n15_w7, 
            w8=> c1_n15_w8, 
            w9=> c1_n15_w9, 
            w10=> c1_n15_w10, 
            w11=> c1_n15_w11, 
            w12=> c1_n15_w12, 
            w13=> c1_n15_w13, 
            w14=> c1_n15_w14, 
            w15=> c1_n15_w15, 
            w16=> c1_n15_w16, 
            w17=> c1_n15_w17, 
            w18=> c1_n15_w18, 
            w19=> c1_n15_w19, 
            w20=> c1_n15_w20, 
            w21=> c1_n15_w21, 
            w22=> c1_n15_w22, 
            w23=> c1_n15_w23, 
            w24=> c1_n15_w24, 
            w25=> c1_n15_w25, 
            w26=> c1_n15_w26, 
            w27=> c1_n15_w27, 
            w28=> c1_n15_w28, 
            w29=> c1_n15_w29, 
            w30=> c1_n15_w30, 
            w31=> c1_n15_w31, 
            w32=> c1_n15_w32, 
            w33=> c1_n15_w33, 
            w34=> c1_n15_w34, 
            w35=> c1_n15_w35, 
            w36=> c1_n15_w36, 
            w37=> c1_n15_w37, 
            w38=> c1_n15_w38, 
            w39=> c1_n15_w39, 
            w40=> c1_n15_w40, 
            w41=> c1_n15_w41, 
            w42=> c1_n15_w42, 
            w43=> c1_n15_w43, 
            w44=> c1_n15_w44, 
            w45=> c1_n15_w45, 
            w46=> c1_n15_w46, 
            w47=> c1_n15_w47, 
            w48=> c1_n15_w48, 
            w49=> c1_n15_w49, 
            w50=> c1_n15_w50, 
            w51=> c1_n15_w51, 
            w52=> c1_n15_w52, 
            w53=> c1_n15_w53, 
            w54=> c1_n15_w54, 
            w55=> c1_n15_w55, 
            w56=> c1_n15_w56, 
            w57=> c1_n15_w57, 
            w58=> c1_n15_w58, 
            w59=> c1_n15_w59, 
            w60=> c1_n15_w60, 
            w61=> c1_n15_w61, 
            w62=> c1_n15_w62, 
            w63=> c1_n15_w63, 
            w64=> c1_n15_w64, 
            w65=> c1_n15_w65, 
            w66=> c1_n15_w66, 
            w67=> c1_n15_w67, 
            w68=> c1_n15_w68, 
            w69=> c1_n15_w69, 
            w70=> c1_n15_w70, 
            w71=> c1_n15_w71, 
            w72=> c1_n15_w72, 
            w73=> c1_n15_w73, 
            w74=> c1_n15_w74, 
            w75=> c1_n15_w75, 
            w76=> c1_n15_w76, 
            w77=> c1_n15_w77, 
            w78=> c1_n15_w78, 
            w79=> c1_n15_w79, 
            w80=> c1_n15_w80, 
            w81=> c1_n15_w81, 
            w82=> c1_n15_w82, 
            w83=> c1_n15_w83, 
            w84=> c1_n15_w84, 
            w85=> c1_n15_w85, 
            w86=> c1_n15_w86, 
            w87=> c1_n15_w87, 
            w88=> c1_n15_w88, 
            w89=> c1_n15_w89, 
            w90=> c1_n15_w90, 
            w91=> c1_n15_w91, 
            w92=> c1_n15_w92, 
            w93=> c1_n15_w93, 
            w94=> c1_n15_w94, 
            w95=> c1_n15_w95, 
            w96=> c1_n15_w96, 
            w97=> c1_n15_w97, 
            w98=> c1_n15_w98, 
            w99=> c1_n15_w99, 
            w100=> c1_n15_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n15_y
   );           
            
neuron_inst_16: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n16_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n16_w1, 
            w2=> c1_n16_w2, 
            w3=> c1_n16_w3, 
            w4=> c1_n16_w4, 
            w5=> c1_n16_w5, 
            w6=> c1_n16_w6, 
            w7=> c1_n16_w7, 
            w8=> c1_n16_w8, 
            w9=> c1_n16_w9, 
            w10=> c1_n16_w10, 
            w11=> c1_n16_w11, 
            w12=> c1_n16_w12, 
            w13=> c1_n16_w13, 
            w14=> c1_n16_w14, 
            w15=> c1_n16_w15, 
            w16=> c1_n16_w16, 
            w17=> c1_n16_w17, 
            w18=> c1_n16_w18, 
            w19=> c1_n16_w19, 
            w20=> c1_n16_w20, 
            w21=> c1_n16_w21, 
            w22=> c1_n16_w22, 
            w23=> c1_n16_w23, 
            w24=> c1_n16_w24, 
            w25=> c1_n16_w25, 
            w26=> c1_n16_w26, 
            w27=> c1_n16_w27, 
            w28=> c1_n16_w28, 
            w29=> c1_n16_w29, 
            w30=> c1_n16_w30, 
            w31=> c1_n16_w31, 
            w32=> c1_n16_w32, 
            w33=> c1_n16_w33, 
            w34=> c1_n16_w34, 
            w35=> c1_n16_w35, 
            w36=> c1_n16_w36, 
            w37=> c1_n16_w37, 
            w38=> c1_n16_w38, 
            w39=> c1_n16_w39, 
            w40=> c1_n16_w40, 
            w41=> c1_n16_w41, 
            w42=> c1_n16_w42, 
            w43=> c1_n16_w43, 
            w44=> c1_n16_w44, 
            w45=> c1_n16_w45, 
            w46=> c1_n16_w46, 
            w47=> c1_n16_w47, 
            w48=> c1_n16_w48, 
            w49=> c1_n16_w49, 
            w50=> c1_n16_w50, 
            w51=> c1_n16_w51, 
            w52=> c1_n16_w52, 
            w53=> c1_n16_w53, 
            w54=> c1_n16_w54, 
            w55=> c1_n16_w55, 
            w56=> c1_n16_w56, 
            w57=> c1_n16_w57, 
            w58=> c1_n16_w58, 
            w59=> c1_n16_w59, 
            w60=> c1_n16_w60, 
            w61=> c1_n16_w61, 
            w62=> c1_n16_w62, 
            w63=> c1_n16_w63, 
            w64=> c1_n16_w64, 
            w65=> c1_n16_w65, 
            w66=> c1_n16_w66, 
            w67=> c1_n16_w67, 
            w68=> c1_n16_w68, 
            w69=> c1_n16_w69, 
            w70=> c1_n16_w70, 
            w71=> c1_n16_w71, 
            w72=> c1_n16_w72, 
            w73=> c1_n16_w73, 
            w74=> c1_n16_w74, 
            w75=> c1_n16_w75, 
            w76=> c1_n16_w76, 
            w77=> c1_n16_w77, 
            w78=> c1_n16_w78, 
            w79=> c1_n16_w79, 
            w80=> c1_n16_w80, 
            w81=> c1_n16_w81, 
            w82=> c1_n16_w82, 
            w83=> c1_n16_w83, 
            w84=> c1_n16_w84, 
            w85=> c1_n16_w85, 
            w86=> c1_n16_w86, 
            w87=> c1_n16_w87, 
            w88=> c1_n16_w88, 
            w89=> c1_n16_w89, 
            w90=> c1_n16_w90, 
            w91=> c1_n16_w91, 
            w92=> c1_n16_w92, 
            w93=> c1_n16_w93, 
            w94=> c1_n16_w94, 
            w95=> c1_n16_w95, 
            w96=> c1_n16_w96, 
            w97=> c1_n16_w97, 
            w98=> c1_n16_w98, 
            w99=> c1_n16_w99, 
            w100=> c1_n16_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n16_y
   );           
            
neuron_inst_17: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n17_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n17_w1, 
            w2=> c1_n17_w2, 
            w3=> c1_n17_w3, 
            w4=> c1_n17_w4, 
            w5=> c1_n17_w5, 
            w6=> c1_n17_w6, 
            w7=> c1_n17_w7, 
            w8=> c1_n17_w8, 
            w9=> c1_n17_w9, 
            w10=> c1_n17_w10, 
            w11=> c1_n17_w11, 
            w12=> c1_n17_w12, 
            w13=> c1_n17_w13, 
            w14=> c1_n17_w14, 
            w15=> c1_n17_w15, 
            w16=> c1_n17_w16, 
            w17=> c1_n17_w17, 
            w18=> c1_n17_w18, 
            w19=> c1_n17_w19, 
            w20=> c1_n17_w20, 
            w21=> c1_n17_w21, 
            w22=> c1_n17_w22, 
            w23=> c1_n17_w23, 
            w24=> c1_n17_w24, 
            w25=> c1_n17_w25, 
            w26=> c1_n17_w26, 
            w27=> c1_n17_w27, 
            w28=> c1_n17_w28, 
            w29=> c1_n17_w29, 
            w30=> c1_n17_w30, 
            w31=> c1_n17_w31, 
            w32=> c1_n17_w32, 
            w33=> c1_n17_w33, 
            w34=> c1_n17_w34, 
            w35=> c1_n17_w35, 
            w36=> c1_n17_w36, 
            w37=> c1_n17_w37, 
            w38=> c1_n17_w38, 
            w39=> c1_n17_w39, 
            w40=> c1_n17_w40, 
            w41=> c1_n17_w41, 
            w42=> c1_n17_w42, 
            w43=> c1_n17_w43, 
            w44=> c1_n17_w44, 
            w45=> c1_n17_w45, 
            w46=> c1_n17_w46, 
            w47=> c1_n17_w47, 
            w48=> c1_n17_w48, 
            w49=> c1_n17_w49, 
            w50=> c1_n17_w50, 
            w51=> c1_n17_w51, 
            w52=> c1_n17_w52, 
            w53=> c1_n17_w53, 
            w54=> c1_n17_w54, 
            w55=> c1_n17_w55, 
            w56=> c1_n17_w56, 
            w57=> c1_n17_w57, 
            w58=> c1_n17_w58, 
            w59=> c1_n17_w59, 
            w60=> c1_n17_w60, 
            w61=> c1_n17_w61, 
            w62=> c1_n17_w62, 
            w63=> c1_n17_w63, 
            w64=> c1_n17_w64, 
            w65=> c1_n17_w65, 
            w66=> c1_n17_w66, 
            w67=> c1_n17_w67, 
            w68=> c1_n17_w68, 
            w69=> c1_n17_w69, 
            w70=> c1_n17_w70, 
            w71=> c1_n17_w71, 
            w72=> c1_n17_w72, 
            w73=> c1_n17_w73, 
            w74=> c1_n17_w74, 
            w75=> c1_n17_w75, 
            w76=> c1_n17_w76, 
            w77=> c1_n17_w77, 
            w78=> c1_n17_w78, 
            w79=> c1_n17_w79, 
            w80=> c1_n17_w80, 
            w81=> c1_n17_w81, 
            w82=> c1_n17_w82, 
            w83=> c1_n17_w83, 
            w84=> c1_n17_w84, 
            w85=> c1_n17_w85, 
            w86=> c1_n17_w86, 
            w87=> c1_n17_w87, 
            w88=> c1_n17_w88, 
            w89=> c1_n17_w89, 
            w90=> c1_n17_w90, 
            w91=> c1_n17_w91, 
            w92=> c1_n17_w92, 
            w93=> c1_n17_w93, 
            w94=> c1_n17_w94, 
            w95=> c1_n17_w95, 
            w96=> c1_n17_w96, 
            w97=> c1_n17_w97, 
            w98=> c1_n17_w98, 
            w99=> c1_n17_w99, 
            w100=> c1_n17_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n17_y
   );           
            
neuron_inst_18: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n18_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n18_w1, 
            w2=> c1_n18_w2, 
            w3=> c1_n18_w3, 
            w4=> c1_n18_w4, 
            w5=> c1_n18_w5, 
            w6=> c1_n18_w6, 
            w7=> c1_n18_w7, 
            w8=> c1_n18_w8, 
            w9=> c1_n18_w9, 
            w10=> c1_n18_w10, 
            w11=> c1_n18_w11, 
            w12=> c1_n18_w12, 
            w13=> c1_n18_w13, 
            w14=> c1_n18_w14, 
            w15=> c1_n18_w15, 
            w16=> c1_n18_w16, 
            w17=> c1_n18_w17, 
            w18=> c1_n18_w18, 
            w19=> c1_n18_w19, 
            w20=> c1_n18_w20, 
            w21=> c1_n18_w21, 
            w22=> c1_n18_w22, 
            w23=> c1_n18_w23, 
            w24=> c1_n18_w24, 
            w25=> c1_n18_w25, 
            w26=> c1_n18_w26, 
            w27=> c1_n18_w27, 
            w28=> c1_n18_w28, 
            w29=> c1_n18_w29, 
            w30=> c1_n18_w30, 
            w31=> c1_n18_w31, 
            w32=> c1_n18_w32, 
            w33=> c1_n18_w33, 
            w34=> c1_n18_w34, 
            w35=> c1_n18_w35, 
            w36=> c1_n18_w36, 
            w37=> c1_n18_w37, 
            w38=> c1_n18_w38, 
            w39=> c1_n18_w39, 
            w40=> c1_n18_w40, 
            w41=> c1_n18_w41, 
            w42=> c1_n18_w42, 
            w43=> c1_n18_w43, 
            w44=> c1_n18_w44, 
            w45=> c1_n18_w45, 
            w46=> c1_n18_w46, 
            w47=> c1_n18_w47, 
            w48=> c1_n18_w48, 
            w49=> c1_n18_w49, 
            w50=> c1_n18_w50, 
            w51=> c1_n18_w51, 
            w52=> c1_n18_w52, 
            w53=> c1_n18_w53, 
            w54=> c1_n18_w54, 
            w55=> c1_n18_w55, 
            w56=> c1_n18_w56, 
            w57=> c1_n18_w57, 
            w58=> c1_n18_w58, 
            w59=> c1_n18_w59, 
            w60=> c1_n18_w60, 
            w61=> c1_n18_w61, 
            w62=> c1_n18_w62, 
            w63=> c1_n18_w63, 
            w64=> c1_n18_w64, 
            w65=> c1_n18_w65, 
            w66=> c1_n18_w66, 
            w67=> c1_n18_w67, 
            w68=> c1_n18_w68, 
            w69=> c1_n18_w69, 
            w70=> c1_n18_w70, 
            w71=> c1_n18_w71, 
            w72=> c1_n18_w72, 
            w73=> c1_n18_w73, 
            w74=> c1_n18_w74, 
            w75=> c1_n18_w75, 
            w76=> c1_n18_w76, 
            w77=> c1_n18_w77, 
            w78=> c1_n18_w78, 
            w79=> c1_n18_w79, 
            w80=> c1_n18_w80, 
            w81=> c1_n18_w81, 
            w82=> c1_n18_w82, 
            w83=> c1_n18_w83, 
            w84=> c1_n18_w84, 
            w85=> c1_n18_w85, 
            w86=> c1_n18_w86, 
            w87=> c1_n18_w87, 
            w88=> c1_n18_w88, 
            w89=> c1_n18_w89, 
            w90=> c1_n18_w90, 
            w91=> c1_n18_w91, 
            w92=> c1_n18_w92, 
            w93=> c1_n18_w93, 
            w94=> c1_n18_w94, 
            w95=> c1_n18_w95, 
            w96=> c1_n18_w96, 
            w97=> c1_n18_w97, 
            w98=> c1_n18_w98, 
            w99=> c1_n18_w99, 
            w100=> c1_n18_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n18_y
   );           
            
neuron_inst_19: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n19_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n19_w1, 
            w2=> c1_n19_w2, 
            w3=> c1_n19_w3, 
            w4=> c1_n19_w4, 
            w5=> c1_n19_w5, 
            w6=> c1_n19_w6, 
            w7=> c1_n19_w7, 
            w8=> c1_n19_w8, 
            w9=> c1_n19_w9, 
            w10=> c1_n19_w10, 
            w11=> c1_n19_w11, 
            w12=> c1_n19_w12, 
            w13=> c1_n19_w13, 
            w14=> c1_n19_w14, 
            w15=> c1_n19_w15, 
            w16=> c1_n19_w16, 
            w17=> c1_n19_w17, 
            w18=> c1_n19_w18, 
            w19=> c1_n19_w19, 
            w20=> c1_n19_w20, 
            w21=> c1_n19_w21, 
            w22=> c1_n19_w22, 
            w23=> c1_n19_w23, 
            w24=> c1_n19_w24, 
            w25=> c1_n19_w25, 
            w26=> c1_n19_w26, 
            w27=> c1_n19_w27, 
            w28=> c1_n19_w28, 
            w29=> c1_n19_w29, 
            w30=> c1_n19_w30, 
            w31=> c1_n19_w31, 
            w32=> c1_n19_w32, 
            w33=> c1_n19_w33, 
            w34=> c1_n19_w34, 
            w35=> c1_n19_w35, 
            w36=> c1_n19_w36, 
            w37=> c1_n19_w37, 
            w38=> c1_n19_w38, 
            w39=> c1_n19_w39, 
            w40=> c1_n19_w40, 
            w41=> c1_n19_w41, 
            w42=> c1_n19_w42, 
            w43=> c1_n19_w43, 
            w44=> c1_n19_w44, 
            w45=> c1_n19_w45, 
            w46=> c1_n19_w46, 
            w47=> c1_n19_w47, 
            w48=> c1_n19_w48, 
            w49=> c1_n19_w49, 
            w50=> c1_n19_w50, 
            w51=> c1_n19_w51, 
            w52=> c1_n19_w52, 
            w53=> c1_n19_w53, 
            w54=> c1_n19_w54, 
            w55=> c1_n19_w55, 
            w56=> c1_n19_w56, 
            w57=> c1_n19_w57, 
            w58=> c1_n19_w58, 
            w59=> c1_n19_w59, 
            w60=> c1_n19_w60, 
            w61=> c1_n19_w61, 
            w62=> c1_n19_w62, 
            w63=> c1_n19_w63, 
            w64=> c1_n19_w64, 
            w65=> c1_n19_w65, 
            w66=> c1_n19_w66, 
            w67=> c1_n19_w67, 
            w68=> c1_n19_w68, 
            w69=> c1_n19_w69, 
            w70=> c1_n19_w70, 
            w71=> c1_n19_w71, 
            w72=> c1_n19_w72, 
            w73=> c1_n19_w73, 
            w74=> c1_n19_w74, 
            w75=> c1_n19_w75, 
            w76=> c1_n19_w76, 
            w77=> c1_n19_w77, 
            w78=> c1_n19_w78, 
            w79=> c1_n19_w79, 
            w80=> c1_n19_w80, 
            w81=> c1_n19_w81, 
            w82=> c1_n19_w82, 
            w83=> c1_n19_w83, 
            w84=> c1_n19_w84, 
            w85=> c1_n19_w85, 
            w86=> c1_n19_w86, 
            w87=> c1_n19_w87, 
            w88=> c1_n19_w88, 
            w89=> c1_n19_w89, 
            w90=> c1_n19_w90, 
            w91=> c1_n19_w91, 
            w92=> c1_n19_w92, 
            w93=> c1_n19_w93, 
            w94=> c1_n19_w94, 
            w95=> c1_n19_w95, 
            w96=> c1_n19_w96, 
            w97=> c1_n19_w97, 
            w98=> c1_n19_w98, 
            w99=> c1_n19_w99, 
            w100=> c1_n19_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n19_y
   );           
            
neuron_inst_20: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n20_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n20_w1, 
            w2=> c1_n20_w2, 
            w3=> c1_n20_w3, 
            w4=> c1_n20_w4, 
            w5=> c1_n20_w5, 
            w6=> c1_n20_w6, 
            w7=> c1_n20_w7, 
            w8=> c1_n20_w8, 
            w9=> c1_n20_w9, 
            w10=> c1_n20_w10, 
            w11=> c1_n20_w11, 
            w12=> c1_n20_w12, 
            w13=> c1_n20_w13, 
            w14=> c1_n20_w14, 
            w15=> c1_n20_w15, 
            w16=> c1_n20_w16, 
            w17=> c1_n20_w17, 
            w18=> c1_n20_w18, 
            w19=> c1_n20_w19, 
            w20=> c1_n20_w20, 
            w21=> c1_n20_w21, 
            w22=> c1_n20_w22, 
            w23=> c1_n20_w23, 
            w24=> c1_n20_w24, 
            w25=> c1_n20_w25, 
            w26=> c1_n20_w26, 
            w27=> c1_n20_w27, 
            w28=> c1_n20_w28, 
            w29=> c1_n20_w29, 
            w30=> c1_n20_w30, 
            w31=> c1_n20_w31, 
            w32=> c1_n20_w32, 
            w33=> c1_n20_w33, 
            w34=> c1_n20_w34, 
            w35=> c1_n20_w35, 
            w36=> c1_n20_w36, 
            w37=> c1_n20_w37, 
            w38=> c1_n20_w38, 
            w39=> c1_n20_w39, 
            w40=> c1_n20_w40, 
            w41=> c1_n20_w41, 
            w42=> c1_n20_w42, 
            w43=> c1_n20_w43, 
            w44=> c1_n20_w44, 
            w45=> c1_n20_w45, 
            w46=> c1_n20_w46, 
            w47=> c1_n20_w47, 
            w48=> c1_n20_w48, 
            w49=> c1_n20_w49, 
            w50=> c1_n20_w50, 
            w51=> c1_n20_w51, 
            w52=> c1_n20_w52, 
            w53=> c1_n20_w53, 
            w54=> c1_n20_w54, 
            w55=> c1_n20_w55, 
            w56=> c1_n20_w56, 
            w57=> c1_n20_w57, 
            w58=> c1_n20_w58, 
            w59=> c1_n20_w59, 
            w60=> c1_n20_w60, 
            w61=> c1_n20_w61, 
            w62=> c1_n20_w62, 
            w63=> c1_n20_w63, 
            w64=> c1_n20_w64, 
            w65=> c1_n20_w65, 
            w66=> c1_n20_w66, 
            w67=> c1_n20_w67, 
            w68=> c1_n20_w68, 
            w69=> c1_n20_w69, 
            w70=> c1_n20_w70, 
            w71=> c1_n20_w71, 
            w72=> c1_n20_w72, 
            w73=> c1_n20_w73, 
            w74=> c1_n20_w74, 
            w75=> c1_n20_w75, 
            w76=> c1_n20_w76, 
            w77=> c1_n20_w77, 
            w78=> c1_n20_w78, 
            w79=> c1_n20_w79, 
            w80=> c1_n20_w80, 
            w81=> c1_n20_w81, 
            w82=> c1_n20_w82, 
            w83=> c1_n20_w83, 
            w84=> c1_n20_w84, 
            w85=> c1_n20_w85, 
            w86=> c1_n20_w86, 
            w87=> c1_n20_w87, 
            w88=> c1_n20_w88, 
            w89=> c1_n20_w89, 
            w90=> c1_n20_w90, 
            w91=> c1_n20_w91, 
            w92=> c1_n20_w92, 
            w93=> c1_n20_w93, 
            w94=> c1_n20_w94, 
            w95=> c1_n20_w95, 
            w96=> c1_n20_w96, 
            w97=> c1_n20_w97, 
            w98=> c1_n20_w98, 
            w99=> c1_n20_w99, 
            w100=> c1_n20_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n20_y
   );           
            
neuron_inst_21: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n21_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n21_w1, 
            w2=> c1_n21_w2, 
            w3=> c1_n21_w3, 
            w4=> c1_n21_w4, 
            w5=> c1_n21_w5, 
            w6=> c1_n21_w6, 
            w7=> c1_n21_w7, 
            w8=> c1_n21_w8, 
            w9=> c1_n21_w9, 
            w10=> c1_n21_w10, 
            w11=> c1_n21_w11, 
            w12=> c1_n21_w12, 
            w13=> c1_n21_w13, 
            w14=> c1_n21_w14, 
            w15=> c1_n21_w15, 
            w16=> c1_n21_w16, 
            w17=> c1_n21_w17, 
            w18=> c1_n21_w18, 
            w19=> c1_n21_w19, 
            w20=> c1_n21_w20, 
            w21=> c1_n21_w21, 
            w22=> c1_n21_w22, 
            w23=> c1_n21_w23, 
            w24=> c1_n21_w24, 
            w25=> c1_n21_w25, 
            w26=> c1_n21_w26, 
            w27=> c1_n21_w27, 
            w28=> c1_n21_w28, 
            w29=> c1_n21_w29, 
            w30=> c1_n21_w30, 
            w31=> c1_n21_w31, 
            w32=> c1_n21_w32, 
            w33=> c1_n21_w33, 
            w34=> c1_n21_w34, 
            w35=> c1_n21_w35, 
            w36=> c1_n21_w36, 
            w37=> c1_n21_w37, 
            w38=> c1_n21_w38, 
            w39=> c1_n21_w39, 
            w40=> c1_n21_w40, 
            w41=> c1_n21_w41, 
            w42=> c1_n21_w42, 
            w43=> c1_n21_w43, 
            w44=> c1_n21_w44, 
            w45=> c1_n21_w45, 
            w46=> c1_n21_w46, 
            w47=> c1_n21_w47, 
            w48=> c1_n21_w48, 
            w49=> c1_n21_w49, 
            w50=> c1_n21_w50, 
            w51=> c1_n21_w51, 
            w52=> c1_n21_w52, 
            w53=> c1_n21_w53, 
            w54=> c1_n21_w54, 
            w55=> c1_n21_w55, 
            w56=> c1_n21_w56, 
            w57=> c1_n21_w57, 
            w58=> c1_n21_w58, 
            w59=> c1_n21_w59, 
            w60=> c1_n21_w60, 
            w61=> c1_n21_w61, 
            w62=> c1_n21_w62, 
            w63=> c1_n21_w63, 
            w64=> c1_n21_w64, 
            w65=> c1_n21_w65, 
            w66=> c1_n21_w66, 
            w67=> c1_n21_w67, 
            w68=> c1_n21_w68, 
            w69=> c1_n21_w69, 
            w70=> c1_n21_w70, 
            w71=> c1_n21_w71, 
            w72=> c1_n21_w72, 
            w73=> c1_n21_w73, 
            w74=> c1_n21_w74, 
            w75=> c1_n21_w75, 
            w76=> c1_n21_w76, 
            w77=> c1_n21_w77, 
            w78=> c1_n21_w78, 
            w79=> c1_n21_w79, 
            w80=> c1_n21_w80, 
            w81=> c1_n21_w81, 
            w82=> c1_n21_w82, 
            w83=> c1_n21_w83, 
            w84=> c1_n21_w84, 
            w85=> c1_n21_w85, 
            w86=> c1_n21_w86, 
            w87=> c1_n21_w87, 
            w88=> c1_n21_w88, 
            w89=> c1_n21_w89, 
            w90=> c1_n21_w90, 
            w91=> c1_n21_w91, 
            w92=> c1_n21_w92, 
            w93=> c1_n21_w93, 
            w94=> c1_n21_w94, 
            w95=> c1_n21_w95, 
            w96=> c1_n21_w96, 
            w97=> c1_n21_w97, 
            w98=> c1_n21_w98, 
            w99=> c1_n21_w99, 
            w100=> c1_n21_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n21_y
   );           
            
neuron_inst_22: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n22_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n22_w1, 
            w2=> c1_n22_w2, 
            w3=> c1_n22_w3, 
            w4=> c1_n22_w4, 
            w5=> c1_n22_w5, 
            w6=> c1_n22_w6, 
            w7=> c1_n22_w7, 
            w8=> c1_n22_w8, 
            w9=> c1_n22_w9, 
            w10=> c1_n22_w10, 
            w11=> c1_n22_w11, 
            w12=> c1_n22_w12, 
            w13=> c1_n22_w13, 
            w14=> c1_n22_w14, 
            w15=> c1_n22_w15, 
            w16=> c1_n22_w16, 
            w17=> c1_n22_w17, 
            w18=> c1_n22_w18, 
            w19=> c1_n22_w19, 
            w20=> c1_n22_w20, 
            w21=> c1_n22_w21, 
            w22=> c1_n22_w22, 
            w23=> c1_n22_w23, 
            w24=> c1_n22_w24, 
            w25=> c1_n22_w25, 
            w26=> c1_n22_w26, 
            w27=> c1_n22_w27, 
            w28=> c1_n22_w28, 
            w29=> c1_n22_w29, 
            w30=> c1_n22_w30, 
            w31=> c1_n22_w31, 
            w32=> c1_n22_w32, 
            w33=> c1_n22_w33, 
            w34=> c1_n22_w34, 
            w35=> c1_n22_w35, 
            w36=> c1_n22_w36, 
            w37=> c1_n22_w37, 
            w38=> c1_n22_w38, 
            w39=> c1_n22_w39, 
            w40=> c1_n22_w40, 
            w41=> c1_n22_w41, 
            w42=> c1_n22_w42, 
            w43=> c1_n22_w43, 
            w44=> c1_n22_w44, 
            w45=> c1_n22_w45, 
            w46=> c1_n22_w46, 
            w47=> c1_n22_w47, 
            w48=> c1_n22_w48, 
            w49=> c1_n22_w49, 
            w50=> c1_n22_w50, 
            w51=> c1_n22_w51, 
            w52=> c1_n22_w52, 
            w53=> c1_n22_w53, 
            w54=> c1_n22_w54, 
            w55=> c1_n22_w55, 
            w56=> c1_n22_w56, 
            w57=> c1_n22_w57, 
            w58=> c1_n22_w58, 
            w59=> c1_n22_w59, 
            w60=> c1_n22_w60, 
            w61=> c1_n22_w61, 
            w62=> c1_n22_w62, 
            w63=> c1_n22_w63, 
            w64=> c1_n22_w64, 
            w65=> c1_n22_w65, 
            w66=> c1_n22_w66, 
            w67=> c1_n22_w67, 
            w68=> c1_n22_w68, 
            w69=> c1_n22_w69, 
            w70=> c1_n22_w70, 
            w71=> c1_n22_w71, 
            w72=> c1_n22_w72, 
            w73=> c1_n22_w73, 
            w74=> c1_n22_w74, 
            w75=> c1_n22_w75, 
            w76=> c1_n22_w76, 
            w77=> c1_n22_w77, 
            w78=> c1_n22_w78, 
            w79=> c1_n22_w79, 
            w80=> c1_n22_w80, 
            w81=> c1_n22_w81, 
            w82=> c1_n22_w82, 
            w83=> c1_n22_w83, 
            w84=> c1_n22_w84, 
            w85=> c1_n22_w85, 
            w86=> c1_n22_w86, 
            w87=> c1_n22_w87, 
            w88=> c1_n22_w88, 
            w89=> c1_n22_w89, 
            w90=> c1_n22_w90, 
            w91=> c1_n22_w91, 
            w92=> c1_n22_w92, 
            w93=> c1_n22_w93, 
            w94=> c1_n22_w94, 
            w95=> c1_n22_w95, 
            w96=> c1_n22_w96, 
            w97=> c1_n22_w97, 
            w98=> c1_n22_w98, 
            w99=> c1_n22_w99, 
            w100=> c1_n22_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n22_y
   );           
            
neuron_inst_23: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n23_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n23_w1, 
            w2=> c1_n23_w2, 
            w3=> c1_n23_w3, 
            w4=> c1_n23_w4, 
            w5=> c1_n23_w5, 
            w6=> c1_n23_w6, 
            w7=> c1_n23_w7, 
            w8=> c1_n23_w8, 
            w9=> c1_n23_w9, 
            w10=> c1_n23_w10, 
            w11=> c1_n23_w11, 
            w12=> c1_n23_w12, 
            w13=> c1_n23_w13, 
            w14=> c1_n23_w14, 
            w15=> c1_n23_w15, 
            w16=> c1_n23_w16, 
            w17=> c1_n23_w17, 
            w18=> c1_n23_w18, 
            w19=> c1_n23_w19, 
            w20=> c1_n23_w20, 
            w21=> c1_n23_w21, 
            w22=> c1_n23_w22, 
            w23=> c1_n23_w23, 
            w24=> c1_n23_w24, 
            w25=> c1_n23_w25, 
            w26=> c1_n23_w26, 
            w27=> c1_n23_w27, 
            w28=> c1_n23_w28, 
            w29=> c1_n23_w29, 
            w30=> c1_n23_w30, 
            w31=> c1_n23_w31, 
            w32=> c1_n23_w32, 
            w33=> c1_n23_w33, 
            w34=> c1_n23_w34, 
            w35=> c1_n23_w35, 
            w36=> c1_n23_w36, 
            w37=> c1_n23_w37, 
            w38=> c1_n23_w38, 
            w39=> c1_n23_w39, 
            w40=> c1_n23_w40, 
            w41=> c1_n23_w41, 
            w42=> c1_n23_w42, 
            w43=> c1_n23_w43, 
            w44=> c1_n23_w44, 
            w45=> c1_n23_w45, 
            w46=> c1_n23_w46, 
            w47=> c1_n23_w47, 
            w48=> c1_n23_w48, 
            w49=> c1_n23_w49, 
            w50=> c1_n23_w50, 
            w51=> c1_n23_w51, 
            w52=> c1_n23_w52, 
            w53=> c1_n23_w53, 
            w54=> c1_n23_w54, 
            w55=> c1_n23_w55, 
            w56=> c1_n23_w56, 
            w57=> c1_n23_w57, 
            w58=> c1_n23_w58, 
            w59=> c1_n23_w59, 
            w60=> c1_n23_w60, 
            w61=> c1_n23_w61, 
            w62=> c1_n23_w62, 
            w63=> c1_n23_w63, 
            w64=> c1_n23_w64, 
            w65=> c1_n23_w65, 
            w66=> c1_n23_w66, 
            w67=> c1_n23_w67, 
            w68=> c1_n23_w68, 
            w69=> c1_n23_w69, 
            w70=> c1_n23_w70, 
            w71=> c1_n23_w71, 
            w72=> c1_n23_w72, 
            w73=> c1_n23_w73, 
            w74=> c1_n23_w74, 
            w75=> c1_n23_w75, 
            w76=> c1_n23_w76, 
            w77=> c1_n23_w77, 
            w78=> c1_n23_w78, 
            w79=> c1_n23_w79, 
            w80=> c1_n23_w80, 
            w81=> c1_n23_w81, 
            w82=> c1_n23_w82, 
            w83=> c1_n23_w83, 
            w84=> c1_n23_w84, 
            w85=> c1_n23_w85, 
            w86=> c1_n23_w86, 
            w87=> c1_n23_w87, 
            w88=> c1_n23_w88, 
            w89=> c1_n23_w89, 
            w90=> c1_n23_w90, 
            w91=> c1_n23_w91, 
            w92=> c1_n23_w92, 
            w93=> c1_n23_w93, 
            w94=> c1_n23_w94, 
            w95=> c1_n23_w95, 
            w96=> c1_n23_w96, 
            w97=> c1_n23_w97, 
            w98=> c1_n23_w98, 
            w99=> c1_n23_w99, 
            w100=> c1_n23_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n23_y
   );           
            
neuron_inst_24: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n24_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n24_w1, 
            w2=> c1_n24_w2, 
            w3=> c1_n24_w3, 
            w4=> c1_n24_w4, 
            w5=> c1_n24_w5, 
            w6=> c1_n24_w6, 
            w7=> c1_n24_w7, 
            w8=> c1_n24_w8, 
            w9=> c1_n24_w9, 
            w10=> c1_n24_w10, 
            w11=> c1_n24_w11, 
            w12=> c1_n24_w12, 
            w13=> c1_n24_w13, 
            w14=> c1_n24_w14, 
            w15=> c1_n24_w15, 
            w16=> c1_n24_w16, 
            w17=> c1_n24_w17, 
            w18=> c1_n24_w18, 
            w19=> c1_n24_w19, 
            w20=> c1_n24_w20, 
            w21=> c1_n24_w21, 
            w22=> c1_n24_w22, 
            w23=> c1_n24_w23, 
            w24=> c1_n24_w24, 
            w25=> c1_n24_w25, 
            w26=> c1_n24_w26, 
            w27=> c1_n24_w27, 
            w28=> c1_n24_w28, 
            w29=> c1_n24_w29, 
            w30=> c1_n24_w30, 
            w31=> c1_n24_w31, 
            w32=> c1_n24_w32, 
            w33=> c1_n24_w33, 
            w34=> c1_n24_w34, 
            w35=> c1_n24_w35, 
            w36=> c1_n24_w36, 
            w37=> c1_n24_w37, 
            w38=> c1_n24_w38, 
            w39=> c1_n24_w39, 
            w40=> c1_n24_w40, 
            w41=> c1_n24_w41, 
            w42=> c1_n24_w42, 
            w43=> c1_n24_w43, 
            w44=> c1_n24_w44, 
            w45=> c1_n24_w45, 
            w46=> c1_n24_w46, 
            w47=> c1_n24_w47, 
            w48=> c1_n24_w48, 
            w49=> c1_n24_w49, 
            w50=> c1_n24_w50, 
            w51=> c1_n24_w51, 
            w52=> c1_n24_w52, 
            w53=> c1_n24_w53, 
            w54=> c1_n24_w54, 
            w55=> c1_n24_w55, 
            w56=> c1_n24_w56, 
            w57=> c1_n24_w57, 
            w58=> c1_n24_w58, 
            w59=> c1_n24_w59, 
            w60=> c1_n24_w60, 
            w61=> c1_n24_w61, 
            w62=> c1_n24_w62, 
            w63=> c1_n24_w63, 
            w64=> c1_n24_w64, 
            w65=> c1_n24_w65, 
            w66=> c1_n24_w66, 
            w67=> c1_n24_w67, 
            w68=> c1_n24_w68, 
            w69=> c1_n24_w69, 
            w70=> c1_n24_w70, 
            w71=> c1_n24_w71, 
            w72=> c1_n24_w72, 
            w73=> c1_n24_w73, 
            w74=> c1_n24_w74, 
            w75=> c1_n24_w75, 
            w76=> c1_n24_w76, 
            w77=> c1_n24_w77, 
            w78=> c1_n24_w78, 
            w79=> c1_n24_w79, 
            w80=> c1_n24_w80, 
            w81=> c1_n24_w81, 
            w82=> c1_n24_w82, 
            w83=> c1_n24_w83, 
            w84=> c1_n24_w84, 
            w85=> c1_n24_w85, 
            w86=> c1_n24_w86, 
            w87=> c1_n24_w87, 
            w88=> c1_n24_w88, 
            w89=> c1_n24_w89, 
            w90=> c1_n24_w90, 
            w91=> c1_n24_w91, 
            w92=> c1_n24_w92, 
            w93=> c1_n24_w93, 
            w94=> c1_n24_w94, 
            w95=> c1_n24_w95, 
            w96=> c1_n24_w96, 
            w97=> c1_n24_w97, 
            w98=> c1_n24_w98, 
            w99=> c1_n24_w99, 
            w100=> c1_n24_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n24_y
   );           
            
neuron_inst_25: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n25_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n25_w1, 
            w2=> c1_n25_w2, 
            w3=> c1_n25_w3, 
            w4=> c1_n25_w4, 
            w5=> c1_n25_w5, 
            w6=> c1_n25_w6, 
            w7=> c1_n25_w7, 
            w8=> c1_n25_w8, 
            w9=> c1_n25_w9, 
            w10=> c1_n25_w10, 
            w11=> c1_n25_w11, 
            w12=> c1_n25_w12, 
            w13=> c1_n25_w13, 
            w14=> c1_n25_w14, 
            w15=> c1_n25_w15, 
            w16=> c1_n25_w16, 
            w17=> c1_n25_w17, 
            w18=> c1_n25_w18, 
            w19=> c1_n25_w19, 
            w20=> c1_n25_w20, 
            w21=> c1_n25_w21, 
            w22=> c1_n25_w22, 
            w23=> c1_n25_w23, 
            w24=> c1_n25_w24, 
            w25=> c1_n25_w25, 
            w26=> c1_n25_w26, 
            w27=> c1_n25_w27, 
            w28=> c1_n25_w28, 
            w29=> c1_n25_w29, 
            w30=> c1_n25_w30, 
            w31=> c1_n25_w31, 
            w32=> c1_n25_w32, 
            w33=> c1_n25_w33, 
            w34=> c1_n25_w34, 
            w35=> c1_n25_w35, 
            w36=> c1_n25_w36, 
            w37=> c1_n25_w37, 
            w38=> c1_n25_w38, 
            w39=> c1_n25_w39, 
            w40=> c1_n25_w40, 
            w41=> c1_n25_w41, 
            w42=> c1_n25_w42, 
            w43=> c1_n25_w43, 
            w44=> c1_n25_w44, 
            w45=> c1_n25_w45, 
            w46=> c1_n25_w46, 
            w47=> c1_n25_w47, 
            w48=> c1_n25_w48, 
            w49=> c1_n25_w49, 
            w50=> c1_n25_w50, 
            w51=> c1_n25_w51, 
            w52=> c1_n25_w52, 
            w53=> c1_n25_w53, 
            w54=> c1_n25_w54, 
            w55=> c1_n25_w55, 
            w56=> c1_n25_w56, 
            w57=> c1_n25_w57, 
            w58=> c1_n25_w58, 
            w59=> c1_n25_w59, 
            w60=> c1_n25_w60, 
            w61=> c1_n25_w61, 
            w62=> c1_n25_w62, 
            w63=> c1_n25_w63, 
            w64=> c1_n25_w64, 
            w65=> c1_n25_w65, 
            w66=> c1_n25_w66, 
            w67=> c1_n25_w67, 
            w68=> c1_n25_w68, 
            w69=> c1_n25_w69, 
            w70=> c1_n25_w70, 
            w71=> c1_n25_w71, 
            w72=> c1_n25_w72, 
            w73=> c1_n25_w73, 
            w74=> c1_n25_w74, 
            w75=> c1_n25_w75, 
            w76=> c1_n25_w76, 
            w77=> c1_n25_w77, 
            w78=> c1_n25_w78, 
            w79=> c1_n25_w79, 
            w80=> c1_n25_w80, 
            w81=> c1_n25_w81, 
            w82=> c1_n25_w82, 
            w83=> c1_n25_w83, 
            w84=> c1_n25_w84, 
            w85=> c1_n25_w85, 
            w86=> c1_n25_w86, 
            w87=> c1_n25_w87, 
            w88=> c1_n25_w88, 
            w89=> c1_n25_w89, 
            w90=> c1_n25_w90, 
            w91=> c1_n25_w91, 
            w92=> c1_n25_w92, 
            w93=> c1_n25_w93, 
            w94=> c1_n25_w94, 
            w95=> c1_n25_w95, 
            w96=> c1_n25_w96, 
            w97=> c1_n25_w97, 
            w98=> c1_n25_w98, 
            w99=> c1_n25_w99, 
            w100=> c1_n25_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n25_y
   );           
            
neuron_inst_26: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n26_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n26_w1, 
            w2=> c1_n26_w2, 
            w3=> c1_n26_w3, 
            w4=> c1_n26_w4, 
            w5=> c1_n26_w5, 
            w6=> c1_n26_w6, 
            w7=> c1_n26_w7, 
            w8=> c1_n26_w8, 
            w9=> c1_n26_w9, 
            w10=> c1_n26_w10, 
            w11=> c1_n26_w11, 
            w12=> c1_n26_w12, 
            w13=> c1_n26_w13, 
            w14=> c1_n26_w14, 
            w15=> c1_n26_w15, 
            w16=> c1_n26_w16, 
            w17=> c1_n26_w17, 
            w18=> c1_n26_w18, 
            w19=> c1_n26_w19, 
            w20=> c1_n26_w20, 
            w21=> c1_n26_w21, 
            w22=> c1_n26_w22, 
            w23=> c1_n26_w23, 
            w24=> c1_n26_w24, 
            w25=> c1_n26_w25, 
            w26=> c1_n26_w26, 
            w27=> c1_n26_w27, 
            w28=> c1_n26_w28, 
            w29=> c1_n26_w29, 
            w30=> c1_n26_w30, 
            w31=> c1_n26_w31, 
            w32=> c1_n26_w32, 
            w33=> c1_n26_w33, 
            w34=> c1_n26_w34, 
            w35=> c1_n26_w35, 
            w36=> c1_n26_w36, 
            w37=> c1_n26_w37, 
            w38=> c1_n26_w38, 
            w39=> c1_n26_w39, 
            w40=> c1_n26_w40, 
            w41=> c1_n26_w41, 
            w42=> c1_n26_w42, 
            w43=> c1_n26_w43, 
            w44=> c1_n26_w44, 
            w45=> c1_n26_w45, 
            w46=> c1_n26_w46, 
            w47=> c1_n26_w47, 
            w48=> c1_n26_w48, 
            w49=> c1_n26_w49, 
            w50=> c1_n26_w50, 
            w51=> c1_n26_w51, 
            w52=> c1_n26_w52, 
            w53=> c1_n26_w53, 
            w54=> c1_n26_w54, 
            w55=> c1_n26_w55, 
            w56=> c1_n26_w56, 
            w57=> c1_n26_w57, 
            w58=> c1_n26_w58, 
            w59=> c1_n26_w59, 
            w60=> c1_n26_w60, 
            w61=> c1_n26_w61, 
            w62=> c1_n26_w62, 
            w63=> c1_n26_w63, 
            w64=> c1_n26_w64, 
            w65=> c1_n26_w65, 
            w66=> c1_n26_w66, 
            w67=> c1_n26_w67, 
            w68=> c1_n26_w68, 
            w69=> c1_n26_w69, 
            w70=> c1_n26_w70, 
            w71=> c1_n26_w71, 
            w72=> c1_n26_w72, 
            w73=> c1_n26_w73, 
            w74=> c1_n26_w74, 
            w75=> c1_n26_w75, 
            w76=> c1_n26_w76, 
            w77=> c1_n26_w77, 
            w78=> c1_n26_w78, 
            w79=> c1_n26_w79, 
            w80=> c1_n26_w80, 
            w81=> c1_n26_w81, 
            w82=> c1_n26_w82, 
            w83=> c1_n26_w83, 
            w84=> c1_n26_w84, 
            w85=> c1_n26_w85, 
            w86=> c1_n26_w86, 
            w87=> c1_n26_w87, 
            w88=> c1_n26_w88, 
            w89=> c1_n26_w89, 
            w90=> c1_n26_w90, 
            w91=> c1_n26_w91, 
            w92=> c1_n26_w92, 
            w93=> c1_n26_w93, 
            w94=> c1_n26_w94, 
            w95=> c1_n26_w95, 
            w96=> c1_n26_w96, 
            w97=> c1_n26_w97, 
            w98=> c1_n26_w98, 
            w99=> c1_n26_w99, 
            w100=> c1_n26_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n26_y
   );           
            
neuron_inst_27: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n27_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n27_w1, 
            w2=> c1_n27_w2, 
            w3=> c1_n27_w3, 
            w4=> c1_n27_w4, 
            w5=> c1_n27_w5, 
            w6=> c1_n27_w6, 
            w7=> c1_n27_w7, 
            w8=> c1_n27_w8, 
            w9=> c1_n27_w9, 
            w10=> c1_n27_w10, 
            w11=> c1_n27_w11, 
            w12=> c1_n27_w12, 
            w13=> c1_n27_w13, 
            w14=> c1_n27_w14, 
            w15=> c1_n27_w15, 
            w16=> c1_n27_w16, 
            w17=> c1_n27_w17, 
            w18=> c1_n27_w18, 
            w19=> c1_n27_w19, 
            w20=> c1_n27_w20, 
            w21=> c1_n27_w21, 
            w22=> c1_n27_w22, 
            w23=> c1_n27_w23, 
            w24=> c1_n27_w24, 
            w25=> c1_n27_w25, 
            w26=> c1_n27_w26, 
            w27=> c1_n27_w27, 
            w28=> c1_n27_w28, 
            w29=> c1_n27_w29, 
            w30=> c1_n27_w30, 
            w31=> c1_n27_w31, 
            w32=> c1_n27_w32, 
            w33=> c1_n27_w33, 
            w34=> c1_n27_w34, 
            w35=> c1_n27_w35, 
            w36=> c1_n27_w36, 
            w37=> c1_n27_w37, 
            w38=> c1_n27_w38, 
            w39=> c1_n27_w39, 
            w40=> c1_n27_w40, 
            w41=> c1_n27_w41, 
            w42=> c1_n27_w42, 
            w43=> c1_n27_w43, 
            w44=> c1_n27_w44, 
            w45=> c1_n27_w45, 
            w46=> c1_n27_w46, 
            w47=> c1_n27_w47, 
            w48=> c1_n27_w48, 
            w49=> c1_n27_w49, 
            w50=> c1_n27_w50, 
            w51=> c1_n27_w51, 
            w52=> c1_n27_w52, 
            w53=> c1_n27_w53, 
            w54=> c1_n27_w54, 
            w55=> c1_n27_w55, 
            w56=> c1_n27_w56, 
            w57=> c1_n27_w57, 
            w58=> c1_n27_w58, 
            w59=> c1_n27_w59, 
            w60=> c1_n27_w60, 
            w61=> c1_n27_w61, 
            w62=> c1_n27_w62, 
            w63=> c1_n27_w63, 
            w64=> c1_n27_w64, 
            w65=> c1_n27_w65, 
            w66=> c1_n27_w66, 
            w67=> c1_n27_w67, 
            w68=> c1_n27_w68, 
            w69=> c1_n27_w69, 
            w70=> c1_n27_w70, 
            w71=> c1_n27_w71, 
            w72=> c1_n27_w72, 
            w73=> c1_n27_w73, 
            w74=> c1_n27_w74, 
            w75=> c1_n27_w75, 
            w76=> c1_n27_w76, 
            w77=> c1_n27_w77, 
            w78=> c1_n27_w78, 
            w79=> c1_n27_w79, 
            w80=> c1_n27_w80, 
            w81=> c1_n27_w81, 
            w82=> c1_n27_w82, 
            w83=> c1_n27_w83, 
            w84=> c1_n27_w84, 
            w85=> c1_n27_w85, 
            w86=> c1_n27_w86, 
            w87=> c1_n27_w87, 
            w88=> c1_n27_w88, 
            w89=> c1_n27_w89, 
            w90=> c1_n27_w90, 
            w91=> c1_n27_w91, 
            w92=> c1_n27_w92, 
            w93=> c1_n27_w93, 
            w94=> c1_n27_w94, 
            w95=> c1_n27_w95, 
            w96=> c1_n27_w96, 
            w97=> c1_n27_w97, 
            w98=> c1_n27_w98, 
            w99=> c1_n27_w99, 
            w100=> c1_n27_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n27_y
   );           
            
neuron_inst_28: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n28_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n28_w1, 
            w2=> c1_n28_w2, 
            w3=> c1_n28_w3, 
            w4=> c1_n28_w4, 
            w5=> c1_n28_w5, 
            w6=> c1_n28_w6, 
            w7=> c1_n28_w7, 
            w8=> c1_n28_w8, 
            w9=> c1_n28_w9, 
            w10=> c1_n28_w10, 
            w11=> c1_n28_w11, 
            w12=> c1_n28_w12, 
            w13=> c1_n28_w13, 
            w14=> c1_n28_w14, 
            w15=> c1_n28_w15, 
            w16=> c1_n28_w16, 
            w17=> c1_n28_w17, 
            w18=> c1_n28_w18, 
            w19=> c1_n28_w19, 
            w20=> c1_n28_w20, 
            w21=> c1_n28_w21, 
            w22=> c1_n28_w22, 
            w23=> c1_n28_w23, 
            w24=> c1_n28_w24, 
            w25=> c1_n28_w25, 
            w26=> c1_n28_w26, 
            w27=> c1_n28_w27, 
            w28=> c1_n28_w28, 
            w29=> c1_n28_w29, 
            w30=> c1_n28_w30, 
            w31=> c1_n28_w31, 
            w32=> c1_n28_w32, 
            w33=> c1_n28_w33, 
            w34=> c1_n28_w34, 
            w35=> c1_n28_w35, 
            w36=> c1_n28_w36, 
            w37=> c1_n28_w37, 
            w38=> c1_n28_w38, 
            w39=> c1_n28_w39, 
            w40=> c1_n28_w40, 
            w41=> c1_n28_w41, 
            w42=> c1_n28_w42, 
            w43=> c1_n28_w43, 
            w44=> c1_n28_w44, 
            w45=> c1_n28_w45, 
            w46=> c1_n28_w46, 
            w47=> c1_n28_w47, 
            w48=> c1_n28_w48, 
            w49=> c1_n28_w49, 
            w50=> c1_n28_w50, 
            w51=> c1_n28_w51, 
            w52=> c1_n28_w52, 
            w53=> c1_n28_w53, 
            w54=> c1_n28_w54, 
            w55=> c1_n28_w55, 
            w56=> c1_n28_w56, 
            w57=> c1_n28_w57, 
            w58=> c1_n28_w58, 
            w59=> c1_n28_w59, 
            w60=> c1_n28_w60, 
            w61=> c1_n28_w61, 
            w62=> c1_n28_w62, 
            w63=> c1_n28_w63, 
            w64=> c1_n28_w64, 
            w65=> c1_n28_w65, 
            w66=> c1_n28_w66, 
            w67=> c1_n28_w67, 
            w68=> c1_n28_w68, 
            w69=> c1_n28_w69, 
            w70=> c1_n28_w70, 
            w71=> c1_n28_w71, 
            w72=> c1_n28_w72, 
            w73=> c1_n28_w73, 
            w74=> c1_n28_w74, 
            w75=> c1_n28_w75, 
            w76=> c1_n28_w76, 
            w77=> c1_n28_w77, 
            w78=> c1_n28_w78, 
            w79=> c1_n28_w79, 
            w80=> c1_n28_w80, 
            w81=> c1_n28_w81, 
            w82=> c1_n28_w82, 
            w83=> c1_n28_w83, 
            w84=> c1_n28_w84, 
            w85=> c1_n28_w85, 
            w86=> c1_n28_w86, 
            w87=> c1_n28_w87, 
            w88=> c1_n28_w88, 
            w89=> c1_n28_w89, 
            w90=> c1_n28_w90, 
            w91=> c1_n28_w91, 
            w92=> c1_n28_w92, 
            w93=> c1_n28_w93, 
            w94=> c1_n28_w94, 
            w95=> c1_n28_w95, 
            w96=> c1_n28_w96, 
            w97=> c1_n28_w97, 
            w98=> c1_n28_w98, 
            w99=> c1_n28_w99, 
            w100=> c1_n28_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n28_y
   );           
            
neuron_inst_29: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n29_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n29_w1, 
            w2=> c1_n29_w2, 
            w3=> c1_n29_w3, 
            w4=> c1_n29_w4, 
            w5=> c1_n29_w5, 
            w6=> c1_n29_w6, 
            w7=> c1_n29_w7, 
            w8=> c1_n29_w8, 
            w9=> c1_n29_w9, 
            w10=> c1_n29_w10, 
            w11=> c1_n29_w11, 
            w12=> c1_n29_w12, 
            w13=> c1_n29_w13, 
            w14=> c1_n29_w14, 
            w15=> c1_n29_w15, 
            w16=> c1_n29_w16, 
            w17=> c1_n29_w17, 
            w18=> c1_n29_w18, 
            w19=> c1_n29_w19, 
            w20=> c1_n29_w20, 
            w21=> c1_n29_w21, 
            w22=> c1_n29_w22, 
            w23=> c1_n29_w23, 
            w24=> c1_n29_w24, 
            w25=> c1_n29_w25, 
            w26=> c1_n29_w26, 
            w27=> c1_n29_w27, 
            w28=> c1_n29_w28, 
            w29=> c1_n29_w29, 
            w30=> c1_n29_w30, 
            w31=> c1_n29_w31, 
            w32=> c1_n29_w32, 
            w33=> c1_n29_w33, 
            w34=> c1_n29_w34, 
            w35=> c1_n29_w35, 
            w36=> c1_n29_w36, 
            w37=> c1_n29_w37, 
            w38=> c1_n29_w38, 
            w39=> c1_n29_w39, 
            w40=> c1_n29_w40, 
            w41=> c1_n29_w41, 
            w42=> c1_n29_w42, 
            w43=> c1_n29_w43, 
            w44=> c1_n29_w44, 
            w45=> c1_n29_w45, 
            w46=> c1_n29_w46, 
            w47=> c1_n29_w47, 
            w48=> c1_n29_w48, 
            w49=> c1_n29_w49, 
            w50=> c1_n29_w50, 
            w51=> c1_n29_w51, 
            w52=> c1_n29_w52, 
            w53=> c1_n29_w53, 
            w54=> c1_n29_w54, 
            w55=> c1_n29_w55, 
            w56=> c1_n29_w56, 
            w57=> c1_n29_w57, 
            w58=> c1_n29_w58, 
            w59=> c1_n29_w59, 
            w60=> c1_n29_w60, 
            w61=> c1_n29_w61, 
            w62=> c1_n29_w62, 
            w63=> c1_n29_w63, 
            w64=> c1_n29_w64, 
            w65=> c1_n29_w65, 
            w66=> c1_n29_w66, 
            w67=> c1_n29_w67, 
            w68=> c1_n29_w68, 
            w69=> c1_n29_w69, 
            w70=> c1_n29_w70, 
            w71=> c1_n29_w71, 
            w72=> c1_n29_w72, 
            w73=> c1_n29_w73, 
            w74=> c1_n29_w74, 
            w75=> c1_n29_w75, 
            w76=> c1_n29_w76, 
            w77=> c1_n29_w77, 
            w78=> c1_n29_w78, 
            w79=> c1_n29_w79, 
            w80=> c1_n29_w80, 
            w81=> c1_n29_w81, 
            w82=> c1_n29_w82, 
            w83=> c1_n29_w83, 
            w84=> c1_n29_w84, 
            w85=> c1_n29_w85, 
            w86=> c1_n29_w86, 
            w87=> c1_n29_w87, 
            w88=> c1_n29_w88, 
            w89=> c1_n29_w89, 
            w90=> c1_n29_w90, 
            w91=> c1_n29_w91, 
            w92=> c1_n29_w92, 
            w93=> c1_n29_w93, 
            w94=> c1_n29_w94, 
            w95=> c1_n29_w95, 
            w96=> c1_n29_w96, 
            w97=> c1_n29_w97, 
            w98=> c1_n29_w98, 
            w99=> c1_n29_w99, 
            w100=> c1_n29_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n29_y
   );           
            
neuron_inst_30: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n30_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n30_w1, 
            w2=> c1_n30_w2, 
            w3=> c1_n30_w3, 
            w4=> c1_n30_w4, 
            w5=> c1_n30_w5, 
            w6=> c1_n30_w6, 
            w7=> c1_n30_w7, 
            w8=> c1_n30_w8, 
            w9=> c1_n30_w9, 
            w10=> c1_n30_w10, 
            w11=> c1_n30_w11, 
            w12=> c1_n30_w12, 
            w13=> c1_n30_w13, 
            w14=> c1_n30_w14, 
            w15=> c1_n30_w15, 
            w16=> c1_n30_w16, 
            w17=> c1_n30_w17, 
            w18=> c1_n30_w18, 
            w19=> c1_n30_w19, 
            w20=> c1_n30_w20, 
            w21=> c1_n30_w21, 
            w22=> c1_n30_w22, 
            w23=> c1_n30_w23, 
            w24=> c1_n30_w24, 
            w25=> c1_n30_w25, 
            w26=> c1_n30_w26, 
            w27=> c1_n30_w27, 
            w28=> c1_n30_w28, 
            w29=> c1_n30_w29, 
            w30=> c1_n30_w30, 
            w31=> c1_n30_w31, 
            w32=> c1_n30_w32, 
            w33=> c1_n30_w33, 
            w34=> c1_n30_w34, 
            w35=> c1_n30_w35, 
            w36=> c1_n30_w36, 
            w37=> c1_n30_w37, 
            w38=> c1_n30_w38, 
            w39=> c1_n30_w39, 
            w40=> c1_n30_w40, 
            w41=> c1_n30_w41, 
            w42=> c1_n30_w42, 
            w43=> c1_n30_w43, 
            w44=> c1_n30_w44, 
            w45=> c1_n30_w45, 
            w46=> c1_n30_w46, 
            w47=> c1_n30_w47, 
            w48=> c1_n30_w48, 
            w49=> c1_n30_w49, 
            w50=> c1_n30_w50, 
            w51=> c1_n30_w51, 
            w52=> c1_n30_w52, 
            w53=> c1_n30_w53, 
            w54=> c1_n30_w54, 
            w55=> c1_n30_w55, 
            w56=> c1_n30_w56, 
            w57=> c1_n30_w57, 
            w58=> c1_n30_w58, 
            w59=> c1_n30_w59, 
            w60=> c1_n30_w60, 
            w61=> c1_n30_w61, 
            w62=> c1_n30_w62, 
            w63=> c1_n30_w63, 
            w64=> c1_n30_w64, 
            w65=> c1_n30_w65, 
            w66=> c1_n30_w66, 
            w67=> c1_n30_w67, 
            w68=> c1_n30_w68, 
            w69=> c1_n30_w69, 
            w70=> c1_n30_w70, 
            w71=> c1_n30_w71, 
            w72=> c1_n30_w72, 
            w73=> c1_n30_w73, 
            w74=> c1_n30_w74, 
            w75=> c1_n30_w75, 
            w76=> c1_n30_w76, 
            w77=> c1_n30_w77, 
            w78=> c1_n30_w78, 
            w79=> c1_n30_w79, 
            w80=> c1_n30_w80, 
            w81=> c1_n30_w81, 
            w82=> c1_n30_w82, 
            w83=> c1_n30_w83, 
            w84=> c1_n30_w84, 
            w85=> c1_n30_w85, 
            w86=> c1_n30_w86, 
            w87=> c1_n30_w87, 
            w88=> c1_n30_w88, 
            w89=> c1_n30_w89, 
            w90=> c1_n30_w90, 
            w91=> c1_n30_w91, 
            w92=> c1_n30_w92, 
            w93=> c1_n30_w93, 
            w94=> c1_n30_w94, 
            w95=> c1_n30_w95, 
            w96=> c1_n30_w96, 
            w97=> c1_n30_w97, 
            w98=> c1_n30_w98, 
            w99=> c1_n30_w99, 
            w100=> c1_n30_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n30_y
   );           
            
neuron_inst_31: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n31_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n31_w1, 
            w2=> c1_n31_w2, 
            w3=> c1_n31_w3, 
            w4=> c1_n31_w4, 
            w5=> c1_n31_w5, 
            w6=> c1_n31_w6, 
            w7=> c1_n31_w7, 
            w8=> c1_n31_w8, 
            w9=> c1_n31_w9, 
            w10=> c1_n31_w10, 
            w11=> c1_n31_w11, 
            w12=> c1_n31_w12, 
            w13=> c1_n31_w13, 
            w14=> c1_n31_w14, 
            w15=> c1_n31_w15, 
            w16=> c1_n31_w16, 
            w17=> c1_n31_w17, 
            w18=> c1_n31_w18, 
            w19=> c1_n31_w19, 
            w20=> c1_n31_w20, 
            w21=> c1_n31_w21, 
            w22=> c1_n31_w22, 
            w23=> c1_n31_w23, 
            w24=> c1_n31_w24, 
            w25=> c1_n31_w25, 
            w26=> c1_n31_w26, 
            w27=> c1_n31_w27, 
            w28=> c1_n31_w28, 
            w29=> c1_n31_w29, 
            w30=> c1_n31_w30, 
            w31=> c1_n31_w31, 
            w32=> c1_n31_w32, 
            w33=> c1_n31_w33, 
            w34=> c1_n31_w34, 
            w35=> c1_n31_w35, 
            w36=> c1_n31_w36, 
            w37=> c1_n31_w37, 
            w38=> c1_n31_w38, 
            w39=> c1_n31_w39, 
            w40=> c1_n31_w40, 
            w41=> c1_n31_w41, 
            w42=> c1_n31_w42, 
            w43=> c1_n31_w43, 
            w44=> c1_n31_w44, 
            w45=> c1_n31_w45, 
            w46=> c1_n31_w46, 
            w47=> c1_n31_w47, 
            w48=> c1_n31_w48, 
            w49=> c1_n31_w49, 
            w50=> c1_n31_w50, 
            w51=> c1_n31_w51, 
            w52=> c1_n31_w52, 
            w53=> c1_n31_w53, 
            w54=> c1_n31_w54, 
            w55=> c1_n31_w55, 
            w56=> c1_n31_w56, 
            w57=> c1_n31_w57, 
            w58=> c1_n31_w58, 
            w59=> c1_n31_w59, 
            w60=> c1_n31_w60, 
            w61=> c1_n31_w61, 
            w62=> c1_n31_w62, 
            w63=> c1_n31_w63, 
            w64=> c1_n31_w64, 
            w65=> c1_n31_w65, 
            w66=> c1_n31_w66, 
            w67=> c1_n31_w67, 
            w68=> c1_n31_w68, 
            w69=> c1_n31_w69, 
            w70=> c1_n31_w70, 
            w71=> c1_n31_w71, 
            w72=> c1_n31_w72, 
            w73=> c1_n31_w73, 
            w74=> c1_n31_w74, 
            w75=> c1_n31_w75, 
            w76=> c1_n31_w76, 
            w77=> c1_n31_w77, 
            w78=> c1_n31_w78, 
            w79=> c1_n31_w79, 
            w80=> c1_n31_w80, 
            w81=> c1_n31_w81, 
            w82=> c1_n31_w82, 
            w83=> c1_n31_w83, 
            w84=> c1_n31_w84, 
            w85=> c1_n31_w85, 
            w86=> c1_n31_w86, 
            w87=> c1_n31_w87, 
            w88=> c1_n31_w88, 
            w89=> c1_n31_w89, 
            w90=> c1_n31_w90, 
            w91=> c1_n31_w91, 
            w92=> c1_n31_w92, 
            w93=> c1_n31_w93, 
            w94=> c1_n31_w94, 
            w95=> c1_n31_w95, 
            w96=> c1_n31_w96, 
            w97=> c1_n31_w97, 
            w98=> c1_n31_w98, 
            w99=> c1_n31_w99, 
            w100=> c1_n31_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n31_y
   );           
            
neuron_inst_32: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n32_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n32_w1, 
            w2=> c1_n32_w2, 
            w3=> c1_n32_w3, 
            w4=> c1_n32_w4, 
            w5=> c1_n32_w5, 
            w6=> c1_n32_w6, 
            w7=> c1_n32_w7, 
            w8=> c1_n32_w8, 
            w9=> c1_n32_w9, 
            w10=> c1_n32_w10, 
            w11=> c1_n32_w11, 
            w12=> c1_n32_w12, 
            w13=> c1_n32_w13, 
            w14=> c1_n32_w14, 
            w15=> c1_n32_w15, 
            w16=> c1_n32_w16, 
            w17=> c1_n32_w17, 
            w18=> c1_n32_w18, 
            w19=> c1_n32_w19, 
            w20=> c1_n32_w20, 
            w21=> c1_n32_w21, 
            w22=> c1_n32_w22, 
            w23=> c1_n32_w23, 
            w24=> c1_n32_w24, 
            w25=> c1_n32_w25, 
            w26=> c1_n32_w26, 
            w27=> c1_n32_w27, 
            w28=> c1_n32_w28, 
            w29=> c1_n32_w29, 
            w30=> c1_n32_w30, 
            w31=> c1_n32_w31, 
            w32=> c1_n32_w32, 
            w33=> c1_n32_w33, 
            w34=> c1_n32_w34, 
            w35=> c1_n32_w35, 
            w36=> c1_n32_w36, 
            w37=> c1_n32_w37, 
            w38=> c1_n32_w38, 
            w39=> c1_n32_w39, 
            w40=> c1_n32_w40, 
            w41=> c1_n32_w41, 
            w42=> c1_n32_w42, 
            w43=> c1_n32_w43, 
            w44=> c1_n32_w44, 
            w45=> c1_n32_w45, 
            w46=> c1_n32_w46, 
            w47=> c1_n32_w47, 
            w48=> c1_n32_w48, 
            w49=> c1_n32_w49, 
            w50=> c1_n32_w50, 
            w51=> c1_n32_w51, 
            w52=> c1_n32_w52, 
            w53=> c1_n32_w53, 
            w54=> c1_n32_w54, 
            w55=> c1_n32_w55, 
            w56=> c1_n32_w56, 
            w57=> c1_n32_w57, 
            w58=> c1_n32_w58, 
            w59=> c1_n32_w59, 
            w60=> c1_n32_w60, 
            w61=> c1_n32_w61, 
            w62=> c1_n32_w62, 
            w63=> c1_n32_w63, 
            w64=> c1_n32_w64, 
            w65=> c1_n32_w65, 
            w66=> c1_n32_w66, 
            w67=> c1_n32_w67, 
            w68=> c1_n32_w68, 
            w69=> c1_n32_w69, 
            w70=> c1_n32_w70, 
            w71=> c1_n32_w71, 
            w72=> c1_n32_w72, 
            w73=> c1_n32_w73, 
            w74=> c1_n32_w74, 
            w75=> c1_n32_w75, 
            w76=> c1_n32_w76, 
            w77=> c1_n32_w77, 
            w78=> c1_n32_w78, 
            w79=> c1_n32_w79, 
            w80=> c1_n32_w80, 
            w81=> c1_n32_w81, 
            w82=> c1_n32_w82, 
            w83=> c1_n32_w83, 
            w84=> c1_n32_w84, 
            w85=> c1_n32_w85, 
            w86=> c1_n32_w86, 
            w87=> c1_n32_w87, 
            w88=> c1_n32_w88, 
            w89=> c1_n32_w89, 
            w90=> c1_n32_w90, 
            w91=> c1_n32_w91, 
            w92=> c1_n32_w92, 
            w93=> c1_n32_w93, 
            w94=> c1_n32_w94, 
            w95=> c1_n32_w95, 
            w96=> c1_n32_w96, 
            w97=> c1_n32_w97, 
            w98=> c1_n32_w98, 
            w99=> c1_n32_w99, 
            w100=> c1_n32_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n32_y
   );           
            
neuron_inst_33: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n33_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n33_w1, 
            w2=> c1_n33_w2, 
            w3=> c1_n33_w3, 
            w4=> c1_n33_w4, 
            w5=> c1_n33_w5, 
            w6=> c1_n33_w6, 
            w7=> c1_n33_w7, 
            w8=> c1_n33_w8, 
            w9=> c1_n33_w9, 
            w10=> c1_n33_w10, 
            w11=> c1_n33_w11, 
            w12=> c1_n33_w12, 
            w13=> c1_n33_w13, 
            w14=> c1_n33_w14, 
            w15=> c1_n33_w15, 
            w16=> c1_n33_w16, 
            w17=> c1_n33_w17, 
            w18=> c1_n33_w18, 
            w19=> c1_n33_w19, 
            w20=> c1_n33_w20, 
            w21=> c1_n33_w21, 
            w22=> c1_n33_w22, 
            w23=> c1_n33_w23, 
            w24=> c1_n33_w24, 
            w25=> c1_n33_w25, 
            w26=> c1_n33_w26, 
            w27=> c1_n33_w27, 
            w28=> c1_n33_w28, 
            w29=> c1_n33_w29, 
            w30=> c1_n33_w30, 
            w31=> c1_n33_w31, 
            w32=> c1_n33_w32, 
            w33=> c1_n33_w33, 
            w34=> c1_n33_w34, 
            w35=> c1_n33_w35, 
            w36=> c1_n33_w36, 
            w37=> c1_n33_w37, 
            w38=> c1_n33_w38, 
            w39=> c1_n33_w39, 
            w40=> c1_n33_w40, 
            w41=> c1_n33_w41, 
            w42=> c1_n33_w42, 
            w43=> c1_n33_w43, 
            w44=> c1_n33_w44, 
            w45=> c1_n33_w45, 
            w46=> c1_n33_w46, 
            w47=> c1_n33_w47, 
            w48=> c1_n33_w48, 
            w49=> c1_n33_w49, 
            w50=> c1_n33_w50, 
            w51=> c1_n33_w51, 
            w52=> c1_n33_w52, 
            w53=> c1_n33_w53, 
            w54=> c1_n33_w54, 
            w55=> c1_n33_w55, 
            w56=> c1_n33_w56, 
            w57=> c1_n33_w57, 
            w58=> c1_n33_w58, 
            w59=> c1_n33_w59, 
            w60=> c1_n33_w60, 
            w61=> c1_n33_w61, 
            w62=> c1_n33_w62, 
            w63=> c1_n33_w63, 
            w64=> c1_n33_w64, 
            w65=> c1_n33_w65, 
            w66=> c1_n33_w66, 
            w67=> c1_n33_w67, 
            w68=> c1_n33_w68, 
            w69=> c1_n33_w69, 
            w70=> c1_n33_w70, 
            w71=> c1_n33_w71, 
            w72=> c1_n33_w72, 
            w73=> c1_n33_w73, 
            w74=> c1_n33_w74, 
            w75=> c1_n33_w75, 
            w76=> c1_n33_w76, 
            w77=> c1_n33_w77, 
            w78=> c1_n33_w78, 
            w79=> c1_n33_w79, 
            w80=> c1_n33_w80, 
            w81=> c1_n33_w81, 
            w82=> c1_n33_w82, 
            w83=> c1_n33_w83, 
            w84=> c1_n33_w84, 
            w85=> c1_n33_w85, 
            w86=> c1_n33_w86, 
            w87=> c1_n33_w87, 
            w88=> c1_n33_w88, 
            w89=> c1_n33_w89, 
            w90=> c1_n33_w90, 
            w91=> c1_n33_w91, 
            w92=> c1_n33_w92, 
            w93=> c1_n33_w93, 
            w94=> c1_n33_w94, 
            w95=> c1_n33_w95, 
            w96=> c1_n33_w96, 
            w97=> c1_n33_w97, 
            w98=> c1_n33_w98, 
            w99=> c1_n33_w99, 
            w100=> c1_n33_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n33_y
   );           
            
neuron_inst_34: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n34_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n34_w1, 
            w2=> c1_n34_w2, 
            w3=> c1_n34_w3, 
            w4=> c1_n34_w4, 
            w5=> c1_n34_w5, 
            w6=> c1_n34_w6, 
            w7=> c1_n34_w7, 
            w8=> c1_n34_w8, 
            w9=> c1_n34_w9, 
            w10=> c1_n34_w10, 
            w11=> c1_n34_w11, 
            w12=> c1_n34_w12, 
            w13=> c1_n34_w13, 
            w14=> c1_n34_w14, 
            w15=> c1_n34_w15, 
            w16=> c1_n34_w16, 
            w17=> c1_n34_w17, 
            w18=> c1_n34_w18, 
            w19=> c1_n34_w19, 
            w20=> c1_n34_w20, 
            w21=> c1_n34_w21, 
            w22=> c1_n34_w22, 
            w23=> c1_n34_w23, 
            w24=> c1_n34_w24, 
            w25=> c1_n34_w25, 
            w26=> c1_n34_w26, 
            w27=> c1_n34_w27, 
            w28=> c1_n34_w28, 
            w29=> c1_n34_w29, 
            w30=> c1_n34_w30, 
            w31=> c1_n34_w31, 
            w32=> c1_n34_w32, 
            w33=> c1_n34_w33, 
            w34=> c1_n34_w34, 
            w35=> c1_n34_w35, 
            w36=> c1_n34_w36, 
            w37=> c1_n34_w37, 
            w38=> c1_n34_w38, 
            w39=> c1_n34_w39, 
            w40=> c1_n34_w40, 
            w41=> c1_n34_w41, 
            w42=> c1_n34_w42, 
            w43=> c1_n34_w43, 
            w44=> c1_n34_w44, 
            w45=> c1_n34_w45, 
            w46=> c1_n34_w46, 
            w47=> c1_n34_w47, 
            w48=> c1_n34_w48, 
            w49=> c1_n34_w49, 
            w50=> c1_n34_w50, 
            w51=> c1_n34_w51, 
            w52=> c1_n34_w52, 
            w53=> c1_n34_w53, 
            w54=> c1_n34_w54, 
            w55=> c1_n34_w55, 
            w56=> c1_n34_w56, 
            w57=> c1_n34_w57, 
            w58=> c1_n34_w58, 
            w59=> c1_n34_w59, 
            w60=> c1_n34_w60, 
            w61=> c1_n34_w61, 
            w62=> c1_n34_w62, 
            w63=> c1_n34_w63, 
            w64=> c1_n34_w64, 
            w65=> c1_n34_w65, 
            w66=> c1_n34_w66, 
            w67=> c1_n34_w67, 
            w68=> c1_n34_w68, 
            w69=> c1_n34_w69, 
            w70=> c1_n34_w70, 
            w71=> c1_n34_w71, 
            w72=> c1_n34_w72, 
            w73=> c1_n34_w73, 
            w74=> c1_n34_w74, 
            w75=> c1_n34_w75, 
            w76=> c1_n34_w76, 
            w77=> c1_n34_w77, 
            w78=> c1_n34_w78, 
            w79=> c1_n34_w79, 
            w80=> c1_n34_w80, 
            w81=> c1_n34_w81, 
            w82=> c1_n34_w82, 
            w83=> c1_n34_w83, 
            w84=> c1_n34_w84, 
            w85=> c1_n34_w85, 
            w86=> c1_n34_w86, 
            w87=> c1_n34_w87, 
            w88=> c1_n34_w88, 
            w89=> c1_n34_w89, 
            w90=> c1_n34_w90, 
            w91=> c1_n34_w91, 
            w92=> c1_n34_w92, 
            w93=> c1_n34_w93, 
            w94=> c1_n34_w94, 
            w95=> c1_n34_w95, 
            w96=> c1_n34_w96, 
            w97=> c1_n34_w97, 
            w98=> c1_n34_w98, 
            w99=> c1_n34_w99, 
            w100=> c1_n34_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n34_y
   );           
            
neuron_inst_35: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n35_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n35_w1, 
            w2=> c1_n35_w2, 
            w3=> c1_n35_w3, 
            w4=> c1_n35_w4, 
            w5=> c1_n35_w5, 
            w6=> c1_n35_w6, 
            w7=> c1_n35_w7, 
            w8=> c1_n35_w8, 
            w9=> c1_n35_w9, 
            w10=> c1_n35_w10, 
            w11=> c1_n35_w11, 
            w12=> c1_n35_w12, 
            w13=> c1_n35_w13, 
            w14=> c1_n35_w14, 
            w15=> c1_n35_w15, 
            w16=> c1_n35_w16, 
            w17=> c1_n35_w17, 
            w18=> c1_n35_w18, 
            w19=> c1_n35_w19, 
            w20=> c1_n35_w20, 
            w21=> c1_n35_w21, 
            w22=> c1_n35_w22, 
            w23=> c1_n35_w23, 
            w24=> c1_n35_w24, 
            w25=> c1_n35_w25, 
            w26=> c1_n35_w26, 
            w27=> c1_n35_w27, 
            w28=> c1_n35_w28, 
            w29=> c1_n35_w29, 
            w30=> c1_n35_w30, 
            w31=> c1_n35_w31, 
            w32=> c1_n35_w32, 
            w33=> c1_n35_w33, 
            w34=> c1_n35_w34, 
            w35=> c1_n35_w35, 
            w36=> c1_n35_w36, 
            w37=> c1_n35_w37, 
            w38=> c1_n35_w38, 
            w39=> c1_n35_w39, 
            w40=> c1_n35_w40, 
            w41=> c1_n35_w41, 
            w42=> c1_n35_w42, 
            w43=> c1_n35_w43, 
            w44=> c1_n35_w44, 
            w45=> c1_n35_w45, 
            w46=> c1_n35_w46, 
            w47=> c1_n35_w47, 
            w48=> c1_n35_w48, 
            w49=> c1_n35_w49, 
            w50=> c1_n35_w50, 
            w51=> c1_n35_w51, 
            w52=> c1_n35_w52, 
            w53=> c1_n35_w53, 
            w54=> c1_n35_w54, 
            w55=> c1_n35_w55, 
            w56=> c1_n35_w56, 
            w57=> c1_n35_w57, 
            w58=> c1_n35_w58, 
            w59=> c1_n35_w59, 
            w60=> c1_n35_w60, 
            w61=> c1_n35_w61, 
            w62=> c1_n35_w62, 
            w63=> c1_n35_w63, 
            w64=> c1_n35_w64, 
            w65=> c1_n35_w65, 
            w66=> c1_n35_w66, 
            w67=> c1_n35_w67, 
            w68=> c1_n35_w68, 
            w69=> c1_n35_w69, 
            w70=> c1_n35_w70, 
            w71=> c1_n35_w71, 
            w72=> c1_n35_w72, 
            w73=> c1_n35_w73, 
            w74=> c1_n35_w74, 
            w75=> c1_n35_w75, 
            w76=> c1_n35_w76, 
            w77=> c1_n35_w77, 
            w78=> c1_n35_w78, 
            w79=> c1_n35_w79, 
            w80=> c1_n35_w80, 
            w81=> c1_n35_w81, 
            w82=> c1_n35_w82, 
            w83=> c1_n35_w83, 
            w84=> c1_n35_w84, 
            w85=> c1_n35_w85, 
            w86=> c1_n35_w86, 
            w87=> c1_n35_w87, 
            w88=> c1_n35_w88, 
            w89=> c1_n35_w89, 
            w90=> c1_n35_w90, 
            w91=> c1_n35_w91, 
            w92=> c1_n35_w92, 
            w93=> c1_n35_w93, 
            w94=> c1_n35_w94, 
            w95=> c1_n35_w95, 
            w96=> c1_n35_w96, 
            w97=> c1_n35_w97, 
            w98=> c1_n35_w98, 
            w99=> c1_n35_w99, 
            w100=> c1_n35_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n35_y
   );           
            
neuron_inst_36: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n36_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n36_w1, 
            w2=> c1_n36_w2, 
            w3=> c1_n36_w3, 
            w4=> c1_n36_w4, 
            w5=> c1_n36_w5, 
            w6=> c1_n36_w6, 
            w7=> c1_n36_w7, 
            w8=> c1_n36_w8, 
            w9=> c1_n36_w9, 
            w10=> c1_n36_w10, 
            w11=> c1_n36_w11, 
            w12=> c1_n36_w12, 
            w13=> c1_n36_w13, 
            w14=> c1_n36_w14, 
            w15=> c1_n36_w15, 
            w16=> c1_n36_w16, 
            w17=> c1_n36_w17, 
            w18=> c1_n36_w18, 
            w19=> c1_n36_w19, 
            w20=> c1_n36_w20, 
            w21=> c1_n36_w21, 
            w22=> c1_n36_w22, 
            w23=> c1_n36_w23, 
            w24=> c1_n36_w24, 
            w25=> c1_n36_w25, 
            w26=> c1_n36_w26, 
            w27=> c1_n36_w27, 
            w28=> c1_n36_w28, 
            w29=> c1_n36_w29, 
            w30=> c1_n36_w30, 
            w31=> c1_n36_w31, 
            w32=> c1_n36_w32, 
            w33=> c1_n36_w33, 
            w34=> c1_n36_w34, 
            w35=> c1_n36_w35, 
            w36=> c1_n36_w36, 
            w37=> c1_n36_w37, 
            w38=> c1_n36_w38, 
            w39=> c1_n36_w39, 
            w40=> c1_n36_w40, 
            w41=> c1_n36_w41, 
            w42=> c1_n36_w42, 
            w43=> c1_n36_w43, 
            w44=> c1_n36_w44, 
            w45=> c1_n36_w45, 
            w46=> c1_n36_w46, 
            w47=> c1_n36_w47, 
            w48=> c1_n36_w48, 
            w49=> c1_n36_w49, 
            w50=> c1_n36_w50, 
            w51=> c1_n36_w51, 
            w52=> c1_n36_w52, 
            w53=> c1_n36_w53, 
            w54=> c1_n36_w54, 
            w55=> c1_n36_w55, 
            w56=> c1_n36_w56, 
            w57=> c1_n36_w57, 
            w58=> c1_n36_w58, 
            w59=> c1_n36_w59, 
            w60=> c1_n36_w60, 
            w61=> c1_n36_w61, 
            w62=> c1_n36_w62, 
            w63=> c1_n36_w63, 
            w64=> c1_n36_w64, 
            w65=> c1_n36_w65, 
            w66=> c1_n36_w66, 
            w67=> c1_n36_w67, 
            w68=> c1_n36_w68, 
            w69=> c1_n36_w69, 
            w70=> c1_n36_w70, 
            w71=> c1_n36_w71, 
            w72=> c1_n36_w72, 
            w73=> c1_n36_w73, 
            w74=> c1_n36_w74, 
            w75=> c1_n36_w75, 
            w76=> c1_n36_w76, 
            w77=> c1_n36_w77, 
            w78=> c1_n36_w78, 
            w79=> c1_n36_w79, 
            w80=> c1_n36_w80, 
            w81=> c1_n36_w81, 
            w82=> c1_n36_w82, 
            w83=> c1_n36_w83, 
            w84=> c1_n36_w84, 
            w85=> c1_n36_w85, 
            w86=> c1_n36_w86, 
            w87=> c1_n36_w87, 
            w88=> c1_n36_w88, 
            w89=> c1_n36_w89, 
            w90=> c1_n36_w90, 
            w91=> c1_n36_w91, 
            w92=> c1_n36_w92, 
            w93=> c1_n36_w93, 
            w94=> c1_n36_w94, 
            w95=> c1_n36_w95, 
            w96=> c1_n36_w96, 
            w97=> c1_n36_w97, 
            w98=> c1_n36_w98, 
            w99=> c1_n36_w99, 
            w100=> c1_n36_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n36_y
   );           
            
neuron_inst_37: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n37_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n37_w1, 
            w2=> c1_n37_w2, 
            w3=> c1_n37_w3, 
            w4=> c1_n37_w4, 
            w5=> c1_n37_w5, 
            w6=> c1_n37_w6, 
            w7=> c1_n37_w7, 
            w8=> c1_n37_w8, 
            w9=> c1_n37_w9, 
            w10=> c1_n37_w10, 
            w11=> c1_n37_w11, 
            w12=> c1_n37_w12, 
            w13=> c1_n37_w13, 
            w14=> c1_n37_w14, 
            w15=> c1_n37_w15, 
            w16=> c1_n37_w16, 
            w17=> c1_n37_w17, 
            w18=> c1_n37_w18, 
            w19=> c1_n37_w19, 
            w20=> c1_n37_w20, 
            w21=> c1_n37_w21, 
            w22=> c1_n37_w22, 
            w23=> c1_n37_w23, 
            w24=> c1_n37_w24, 
            w25=> c1_n37_w25, 
            w26=> c1_n37_w26, 
            w27=> c1_n37_w27, 
            w28=> c1_n37_w28, 
            w29=> c1_n37_w29, 
            w30=> c1_n37_w30, 
            w31=> c1_n37_w31, 
            w32=> c1_n37_w32, 
            w33=> c1_n37_w33, 
            w34=> c1_n37_w34, 
            w35=> c1_n37_w35, 
            w36=> c1_n37_w36, 
            w37=> c1_n37_w37, 
            w38=> c1_n37_w38, 
            w39=> c1_n37_w39, 
            w40=> c1_n37_w40, 
            w41=> c1_n37_w41, 
            w42=> c1_n37_w42, 
            w43=> c1_n37_w43, 
            w44=> c1_n37_w44, 
            w45=> c1_n37_w45, 
            w46=> c1_n37_w46, 
            w47=> c1_n37_w47, 
            w48=> c1_n37_w48, 
            w49=> c1_n37_w49, 
            w50=> c1_n37_w50, 
            w51=> c1_n37_w51, 
            w52=> c1_n37_w52, 
            w53=> c1_n37_w53, 
            w54=> c1_n37_w54, 
            w55=> c1_n37_w55, 
            w56=> c1_n37_w56, 
            w57=> c1_n37_w57, 
            w58=> c1_n37_w58, 
            w59=> c1_n37_w59, 
            w60=> c1_n37_w60, 
            w61=> c1_n37_w61, 
            w62=> c1_n37_w62, 
            w63=> c1_n37_w63, 
            w64=> c1_n37_w64, 
            w65=> c1_n37_w65, 
            w66=> c1_n37_w66, 
            w67=> c1_n37_w67, 
            w68=> c1_n37_w68, 
            w69=> c1_n37_w69, 
            w70=> c1_n37_w70, 
            w71=> c1_n37_w71, 
            w72=> c1_n37_w72, 
            w73=> c1_n37_w73, 
            w74=> c1_n37_w74, 
            w75=> c1_n37_w75, 
            w76=> c1_n37_w76, 
            w77=> c1_n37_w77, 
            w78=> c1_n37_w78, 
            w79=> c1_n37_w79, 
            w80=> c1_n37_w80, 
            w81=> c1_n37_w81, 
            w82=> c1_n37_w82, 
            w83=> c1_n37_w83, 
            w84=> c1_n37_w84, 
            w85=> c1_n37_w85, 
            w86=> c1_n37_w86, 
            w87=> c1_n37_w87, 
            w88=> c1_n37_w88, 
            w89=> c1_n37_w89, 
            w90=> c1_n37_w90, 
            w91=> c1_n37_w91, 
            w92=> c1_n37_w92, 
            w93=> c1_n37_w93, 
            w94=> c1_n37_w94, 
            w95=> c1_n37_w95, 
            w96=> c1_n37_w96, 
            w97=> c1_n37_w97, 
            w98=> c1_n37_w98, 
            w99=> c1_n37_w99, 
            w100=> c1_n37_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n37_y
   );           
            
neuron_inst_38: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n38_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n38_w1, 
            w2=> c1_n38_w2, 
            w3=> c1_n38_w3, 
            w4=> c1_n38_w4, 
            w5=> c1_n38_w5, 
            w6=> c1_n38_w6, 
            w7=> c1_n38_w7, 
            w8=> c1_n38_w8, 
            w9=> c1_n38_w9, 
            w10=> c1_n38_w10, 
            w11=> c1_n38_w11, 
            w12=> c1_n38_w12, 
            w13=> c1_n38_w13, 
            w14=> c1_n38_w14, 
            w15=> c1_n38_w15, 
            w16=> c1_n38_w16, 
            w17=> c1_n38_w17, 
            w18=> c1_n38_w18, 
            w19=> c1_n38_w19, 
            w20=> c1_n38_w20, 
            w21=> c1_n38_w21, 
            w22=> c1_n38_w22, 
            w23=> c1_n38_w23, 
            w24=> c1_n38_w24, 
            w25=> c1_n38_w25, 
            w26=> c1_n38_w26, 
            w27=> c1_n38_w27, 
            w28=> c1_n38_w28, 
            w29=> c1_n38_w29, 
            w30=> c1_n38_w30, 
            w31=> c1_n38_w31, 
            w32=> c1_n38_w32, 
            w33=> c1_n38_w33, 
            w34=> c1_n38_w34, 
            w35=> c1_n38_w35, 
            w36=> c1_n38_w36, 
            w37=> c1_n38_w37, 
            w38=> c1_n38_w38, 
            w39=> c1_n38_w39, 
            w40=> c1_n38_w40, 
            w41=> c1_n38_w41, 
            w42=> c1_n38_w42, 
            w43=> c1_n38_w43, 
            w44=> c1_n38_w44, 
            w45=> c1_n38_w45, 
            w46=> c1_n38_w46, 
            w47=> c1_n38_w47, 
            w48=> c1_n38_w48, 
            w49=> c1_n38_w49, 
            w50=> c1_n38_w50, 
            w51=> c1_n38_w51, 
            w52=> c1_n38_w52, 
            w53=> c1_n38_w53, 
            w54=> c1_n38_w54, 
            w55=> c1_n38_w55, 
            w56=> c1_n38_w56, 
            w57=> c1_n38_w57, 
            w58=> c1_n38_w58, 
            w59=> c1_n38_w59, 
            w60=> c1_n38_w60, 
            w61=> c1_n38_w61, 
            w62=> c1_n38_w62, 
            w63=> c1_n38_w63, 
            w64=> c1_n38_w64, 
            w65=> c1_n38_w65, 
            w66=> c1_n38_w66, 
            w67=> c1_n38_w67, 
            w68=> c1_n38_w68, 
            w69=> c1_n38_w69, 
            w70=> c1_n38_w70, 
            w71=> c1_n38_w71, 
            w72=> c1_n38_w72, 
            w73=> c1_n38_w73, 
            w74=> c1_n38_w74, 
            w75=> c1_n38_w75, 
            w76=> c1_n38_w76, 
            w77=> c1_n38_w77, 
            w78=> c1_n38_w78, 
            w79=> c1_n38_w79, 
            w80=> c1_n38_w80, 
            w81=> c1_n38_w81, 
            w82=> c1_n38_w82, 
            w83=> c1_n38_w83, 
            w84=> c1_n38_w84, 
            w85=> c1_n38_w85, 
            w86=> c1_n38_w86, 
            w87=> c1_n38_w87, 
            w88=> c1_n38_w88, 
            w89=> c1_n38_w89, 
            w90=> c1_n38_w90, 
            w91=> c1_n38_w91, 
            w92=> c1_n38_w92, 
            w93=> c1_n38_w93, 
            w94=> c1_n38_w94, 
            w95=> c1_n38_w95, 
            w96=> c1_n38_w96, 
            w97=> c1_n38_w97, 
            w98=> c1_n38_w98, 
            w99=> c1_n38_w99, 
            w100=> c1_n38_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n38_y
   );           
            
neuron_inst_39: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n39_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n39_w1, 
            w2=> c1_n39_w2, 
            w3=> c1_n39_w3, 
            w4=> c1_n39_w4, 
            w5=> c1_n39_w5, 
            w6=> c1_n39_w6, 
            w7=> c1_n39_w7, 
            w8=> c1_n39_w8, 
            w9=> c1_n39_w9, 
            w10=> c1_n39_w10, 
            w11=> c1_n39_w11, 
            w12=> c1_n39_w12, 
            w13=> c1_n39_w13, 
            w14=> c1_n39_w14, 
            w15=> c1_n39_w15, 
            w16=> c1_n39_w16, 
            w17=> c1_n39_w17, 
            w18=> c1_n39_w18, 
            w19=> c1_n39_w19, 
            w20=> c1_n39_w20, 
            w21=> c1_n39_w21, 
            w22=> c1_n39_w22, 
            w23=> c1_n39_w23, 
            w24=> c1_n39_w24, 
            w25=> c1_n39_w25, 
            w26=> c1_n39_w26, 
            w27=> c1_n39_w27, 
            w28=> c1_n39_w28, 
            w29=> c1_n39_w29, 
            w30=> c1_n39_w30, 
            w31=> c1_n39_w31, 
            w32=> c1_n39_w32, 
            w33=> c1_n39_w33, 
            w34=> c1_n39_w34, 
            w35=> c1_n39_w35, 
            w36=> c1_n39_w36, 
            w37=> c1_n39_w37, 
            w38=> c1_n39_w38, 
            w39=> c1_n39_w39, 
            w40=> c1_n39_w40, 
            w41=> c1_n39_w41, 
            w42=> c1_n39_w42, 
            w43=> c1_n39_w43, 
            w44=> c1_n39_w44, 
            w45=> c1_n39_w45, 
            w46=> c1_n39_w46, 
            w47=> c1_n39_w47, 
            w48=> c1_n39_w48, 
            w49=> c1_n39_w49, 
            w50=> c1_n39_w50, 
            w51=> c1_n39_w51, 
            w52=> c1_n39_w52, 
            w53=> c1_n39_w53, 
            w54=> c1_n39_w54, 
            w55=> c1_n39_w55, 
            w56=> c1_n39_w56, 
            w57=> c1_n39_w57, 
            w58=> c1_n39_w58, 
            w59=> c1_n39_w59, 
            w60=> c1_n39_w60, 
            w61=> c1_n39_w61, 
            w62=> c1_n39_w62, 
            w63=> c1_n39_w63, 
            w64=> c1_n39_w64, 
            w65=> c1_n39_w65, 
            w66=> c1_n39_w66, 
            w67=> c1_n39_w67, 
            w68=> c1_n39_w68, 
            w69=> c1_n39_w69, 
            w70=> c1_n39_w70, 
            w71=> c1_n39_w71, 
            w72=> c1_n39_w72, 
            w73=> c1_n39_w73, 
            w74=> c1_n39_w74, 
            w75=> c1_n39_w75, 
            w76=> c1_n39_w76, 
            w77=> c1_n39_w77, 
            w78=> c1_n39_w78, 
            w79=> c1_n39_w79, 
            w80=> c1_n39_w80, 
            w81=> c1_n39_w81, 
            w82=> c1_n39_w82, 
            w83=> c1_n39_w83, 
            w84=> c1_n39_w84, 
            w85=> c1_n39_w85, 
            w86=> c1_n39_w86, 
            w87=> c1_n39_w87, 
            w88=> c1_n39_w88, 
            w89=> c1_n39_w89, 
            w90=> c1_n39_w90, 
            w91=> c1_n39_w91, 
            w92=> c1_n39_w92, 
            w93=> c1_n39_w93, 
            w94=> c1_n39_w94, 
            w95=> c1_n39_w95, 
            w96=> c1_n39_w96, 
            w97=> c1_n39_w97, 
            w98=> c1_n39_w98, 
            w99=> c1_n39_w99, 
            w100=> c1_n39_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n39_y
   );           
            
neuron_inst_40: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n40_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n40_w1, 
            w2=> c1_n40_w2, 
            w3=> c1_n40_w3, 
            w4=> c1_n40_w4, 
            w5=> c1_n40_w5, 
            w6=> c1_n40_w6, 
            w7=> c1_n40_w7, 
            w8=> c1_n40_w8, 
            w9=> c1_n40_w9, 
            w10=> c1_n40_w10, 
            w11=> c1_n40_w11, 
            w12=> c1_n40_w12, 
            w13=> c1_n40_w13, 
            w14=> c1_n40_w14, 
            w15=> c1_n40_w15, 
            w16=> c1_n40_w16, 
            w17=> c1_n40_w17, 
            w18=> c1_n40_w18, 
            w19=> c1_n40_w19, 
            w20=> c1_n40_w20, 
            w21=> c1_n40_w21, 
            w22=> c1_n40_w22, 
            w23=> c1_n40_w23, 
            w24=> c1_n40_w24, 
            w25=> c1_n40_w25, 
            w26=> c1_n40_w26, 
            w27=> c1_n40_w27, 
            w28=> c1_n40_w28, 
            w29=> c1_n40_w29, 
            w30=> c1_n40_w30, 
            w31=> c1_n40_w31, 
            w32=> c1_n40_w32, 
            w33=> c1_n40_w33, 
            w34=> c1_n40_w34, 
            w35=> c1_n40_w35, 
            w36=> c1_n40_w36, 
            w37=> c1_n40_w37, 
            w38=> c1_n40_w38, 
            w39=> c1_n40_w39, 
            w40=> c1_n40_w40, 
            w41=> c1_n40_w41, 
            w42=> c1_n40_w42, 
            w43=> c1_n40_w43, 
            w44=> c1_n40_w44, 
            w45=> c1_n40_w45, 
            w46=> c1_n40_w46, 
            w47=> c1_n40_w47, 
            w48=> c1_n40_w48, 
            w49=> c1_n40_w49, 
            w50=> c1_n40_w50, 
            w51=> c1_n40_w51, 
            w52=> c1_n40_w52, 
            w53=> c1_n40_w53, 
            w54=> c1_n40_w54, 
            w55=> c1_n40_w55, 
            w56=> c1_n40_w56, 
            w57=> c1_n40_w57, 
            w58=> c1_n40_w58, 
            w59=> c1_n40_w59, 
            w60=> c1_n40_w60, 
            w61=> c1_n40_w61, 
            w62=> c1_n40_w62, 
            w63=> c1_n40_w63, 
            w64=> c1_n40_w64, 
            w65=> c1_n40_w65, 
            w66=> c1_n40_w66, 
            w67=> c1_n40_w67, 
            w68=> c1_n40_w68, 
            w69=> c1_n40_w69, 
            w70=> c1_n40_w70, 
            w71=> c1_n40_w71, 
            w72=> c1_n40_w72, 
            w73=> c1_n40_w73, 
            w74=> c1_n40_w74, 
            w75=> c1_n40_w75, 
            w76=> c1_n40_w76, 
            w77=> c1_n40_w77, 
            w78=> c1_n40_w78, 
            w79=> c1_n40_w79, 
            w80=> c1_n40_w80, 
            w81=> c1_n40_w81, 
            w82=> c1_n40_w82, 
            w83=> c1_n40_w83, 
            w84=> c1_n40_w84, 
            w85=> c1_n40_w85, 
            w86=> c1_n40_w86, 
            w87=> c1_n40_w87, 
            w88=> c1_n40_w88, 
            w89=> c1_n40_w89, 
            w90=> c1_n40_w90, 
            w91=> c1_n40_w91, 
            w92=> c1_n40_w92, 
            w93=> c1_n40_w93, 
            w94=> c1_n40_w94, 
            w95=> c1_n40_w95, 
            w96=> c1_n40_w96, 
            w97=> c1_n40_w97, 
            w98=> c1_n40_w98, 
            w99=> c1_n40_w99, 
            w100=> c1_n40_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n40_y
   );           
            
neuron_inst_41: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n41_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n41_w1, 
            w2=> c1_n41_w2, 
            w3=> c1_n41_w3, 
            w4=> c1_n41_w4, 
            w5=> c1_n41_w5, 
            w6=> c1_n41_w6, 
            w7=> c1_n41_w7, 
            w8=> c1_n41_w8, 
            w9=> c1_n41_w9, 
            w10=> c1_n41_w10, 
            w11=> c1_n41_w11, 
            w12=> c1_n41_w12, 
            w13=> c1_n41_w13, 
            w14=> c1_n41_w14, 
            w15=> c1_n41_w15, 
            w16=> c1_n41_w16, 
            w17=> c1_n41_w17, 
            w18=> c1_n41_w18, 
            w19=> c1_n41_w19, 
            w20=> c1_n41_w20, 
            w21=> c1_n41_w21, 
            w22=> c1_n41_w22, 
            w23=> c1_n41_w23, 
            w24=> c1_n41_w24, 
            w25=> c1_n41_w25, 
            w26=> c1_n41_w26, 
            w27=> c1_n41_w27, 
            w28=> c1_n41_w28, 
            w29=> c1_n41_w29, 
            w30=> c1_n41_w30, 
            w31=> c1_n41_w31, 
            w32=> c1_n41_w32, 
            w33=> c1_n41_w33, 
            w34=> c1_n41_w34, 
            w35=> c1_n41_w35, 
            w36=> c1_n41_w36, 
            w37=> c1_n41_w37, 
            w38=> c1_n41_w38, 
            w39=> c1_n41_w39, 
            w40=> c1_n41_w40, 
            w41=> c1_n41_w41, 
            w42=> c1_n41_w42, 
            w43=> c1_n41_w43, 
            w44=> c1_n41_w44, 
            w45=> c1_n41_w45, 
            w46=> c1_n41_w46, 
            w47=> c1_n41_w47, 
            w48=> c1_n41_w48, 
            w49=> c1_n41_w49, 
            w50=> c1_n41_w50, 
            w51=> c1_n41_w51, 
            w52=> c1_n41_w52, 
            w53=> c1_n41_w53, 
            w54=> c1_n41_w54, 
            w55=> c1_n41_w55, 
            w56=> c1_n41_w56, 
            w57=> c1_n41_w57, 
            w58=> c1_n41_w58, 
            w59=> c1_n41_w59, 
            w60=> c1_n41_w60, 
            w61=> c1_n41_w61, 
            w62=> c1_n41_w62, 
            w63=> c1_n41_w63, 
            w64=> c1_n41_w64, 
            w65=> c1_n41_w65, 
            w66=> c1_n41_w66, 
            w67=> c1_n41_w67, 
            w68=> c1_n41_w68, 
            w69=> c1_n41_w69, 
            w70=> c1_n41_w70, 
            w71=> c1_n41_w71, 
            w72=> c1_n41_w72, 
            w73=> c1_n41_w73, 
            w74=> c1_n41_w74, 
            w75=> c1_n41_w75, 
            w76=> c1_n41_w76, 
            w77=> c1_n41_w77, 
            w78=> c1_n41_w78, 
            w79=> c1_n41_w79, 
            w80=> c1_n41_w80, 
            w81=> c1_n41_w81, 
            w82=> c1_n41_w82, 
            w83=> c1_n41_w83, 
            w84=> c1_n41_w84, 
            w85=> c1_n41_w85, 
            w86=> c1_n41_w86, 
            w87=> c1_n41_w87, 
            w88=> c1_n41_w88, 
            w89=> c1_n41_w89, 
            w90=> c1_n41_w90, 
            w91=> c1_n41_w91, 
            w92=> c1_n41_w92, 
            w93=> c1_n41_w93, 
            w94=> c1_n41_w94, 
            w95=> c1_n41_w95, 
            w96=> c1_n41_w96, 
            w97=> c1_n41_w97, 
            w98=> c1_n41_w98, 
            w99=> c1_n41_w99, 
            w100=> c1_n41_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n41_y
   );           
            
neuron_inst_42: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n42_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n42_w1, 
            w2=> c1_n42_w2, 
            w3=> c1_n42_w3, 
            w4=> c1_n42_w4, 
            w5=> c1_n42_w5, 
            w6=> c1_n42_w6, 
            w7=> c1_n42_w7, 
            w8=> c1_n42_w8, 
            w9=> c1_n42_w9, 
            w10=> c1_n42_w10, 
            w11=> c1_n42_w11, 
            w12=> c1_n42_w12, 
            w13=> c1_n42_w13, 
            w14=> c1_n42_w14, 
            w15=> c1_n42_w15, 
            w16=> c1_n42_w16, 
            w17=> c1_n42_w17, 
            w18=> c1_n42_w18, 
            w19=> c1_n42_w19, 
            w20=> c1_n42_w20, 
            w21=> c1_n42_w21, 
            w22=> c1_n42_w22, 
            w23=> c1_n42_w23, 
            w24=> c1_n42_w24, 
            w25=> c1_n42_w25, 
            w26=> c1_n42_w26, 
            w27=> c1_n42_w27, 
            w28=> c1_n42_w28, 
            w29=> c1_n42_w29, 
            w30=> c1_n42_w30, 
            w31=> c1_n42_w31, 
            w32=> c1_n42_w32, 
            w33=> c1_n42_w33, 
            w34=> c1_n42_w34, 
            w35=> c1_n42_w35, 
            w36=> c1_n42_w36, 
            w37=> c1_n42_w37, 
            w38=> c1_n42_w38, 
            w39=> c1_n42_w39, 
            w40=> c1_n42_w40, 
            w41=> c1_n42_w41, 
            w42=> c1_n42_w42, 
            w43=> c1_n42_w43, 
            w44=> c1_n42_w44, 
            w45=> c1_n42_w45, 
            w46=> c1_n42_w46, 
            w47=> c1_n42_w47, 
            w48=> c1_n42_w48, 
            w49=> c1_n42_w49, 
            w50=> c1_n42_w50, 
            w51=> c1_n42_w51, 
            w52=> c1_n42_w52, 
            w53=> c1_n42_w53, 
            w54=> c1_n42_w54, 
            w55=> c1_n42_w55, 
            w56=> c1_n42_w56, 
            w57=> c1_n42_w57, 
            w58=> c1_n42_w58, 
            w59=> c1_n42_w59, 
            w60=> c1_n42_w60, 
            w61=> c1_n42_w61, 
            w62=> c1_n42_w62, 
            w63=> c1_n42_w63, 
            w64=> c1_n42_w64, 
            w65=> c1_n42_w65, 
            w66=> c1_n42_w66, 
            w67=> c1_n42_w67, 
            w68=> c1_n42_w68, 
            w69=> c1_n42_w69, 
            w70=> c1_n42_w70, 
            w71=> c1_n42_w71, 
            w72=> c1_n42_w72, 
            w73=> c1_n42_w73, 
            w74=> c1_n42_w74, 
            w75=> c1_n42_w75, 
            w76=> c1_n42_w76, 
            w77=> c1_n42_w77, 
            w78=> c1_n42_w78, 
            w79=> c1_n42_w79, 
            w80=> c1_n42_w80, 
            w81=> c1_n42_w81, 
            w82=> c1_n42_w82, 
            w83=> c1_n42_w83, 
            w84=> c1_n42_w84, 
            w85=> c1_n42_w85, 
            w86=> c1_n42_w86, 
            w87=> c1_n42_w87, 
            w88=> c1_n42_w88, 
            w89=> c1_n42_w89, 
            w90=> c1_n42_w90, 
            w91=> c1_n42_w91, 
            w92=> c1_n42_w92, 
            w93=> c1_n42_w93, 
            w94=> c1_n42_w94, 
            w95=> c1_n42_w95, 
            w96=> c1_n42_w96, 
            w97=> c1_n42_w97, 
            w98=> c1_n42_w98, 
            w99=> c1_n42_w99, 
            w100=> c1_n42_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n42_y
   );           
            
neuron_inst_43: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n43_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n43_w1, 
            w2=> c1_n43_w2, 
            w3=> c1_n43_w3, 
            w4=> c1_n43_w4, 
            w5=> c1_n43_w5, 
            w6=> c1_n43_w6, 
            w7=> c1_n43_w7, 
            w8=> c1_n43_w8, 
            w9=> c1_n43_w9, 
            w10=> c1_n43_w10, 
            w11=> c1_n43_w11, 
            w12=> c1_n43_w12, 
            w13=> c1_n43_w13, 
            w14=> c1_n43_w14, 
            w15=> c1_n43_w15, 
            w16=> c1_n43_w16, 
            w17=> c1_n43_w17, 
            w18=> c1_n43_w18, 
            w19=> c1_n43_w19, 
            w20=> c1_n43_w20, 
            w21=> c1_n43_w21, 
            w22=> c1_n43_w22, 
            w23=> c1_n43_w23, 
            w24=> c1_n43_w24, 
            w25=> c1_n43_w25, 
            w26=> c1_n43_w26, 
            w27=> c1_n43_w27, 
            w28=> c1_n43_w28, 
            w29=> c1_n43_w29, 
            w30=> c1_n43_w30, 
            w31=> c1_n43_w31, 
            w32=> c1_n43_w32, 
            w33=> c1_n43_w33, 
            w34=> c1_n43_w34, 
            w35=> c1_n43_w35, 
            w36=> c1_n43_w36, 
            w37=> c1_n43_w37, 
            w38=> c1_n43_w38, 
            w39=> c1_n43_w39, 
            w40=> c1_n43_w40, 
            w41=> c1_n43_w41, 
            w42=> c1_n43_w42, 
            w43=> c1_n43_w43, 
            w44=> c1_n43_w44, 
            w45=> c1_n43_w45, 
            w46=> c1_n43_w46, 
            w47=> c1_n43_w47, 
            w48=> c1_n43_w48, 
            w49=> c1_n43_w49, 
            w50=> c1_n43_w50, 
            w51=> c1_n43_w51, 
            w52=> c1_n43_w52, 
            w53=> c1_n43_w53, 
            w54=> c1_n43_w54, 
            w55=> c1_n43_w55, 
            w56=> c1_n43_w56, 
            w57=> c1_n43_w57, 
            w58=> c1_n43_w58, 
            w59=> c1_n43_w59, 
            w60=> c1_n43_w60, 
            w61=> c1_n43_w61, 
            w62=> c1_n43_w62, 
            w63=> c1_n43_w63, 
            w64=> c1_n43_w64, 
            w65=> c1_n43_w65, 
            w66=> c1_n43_w66, 
            w67=> c1_n43_w67, 
            w68=> c1_n43_w68, 
            w69=> c1_n43_w69, 
            w70=> c1_n43_w70, 
            w71=> c1_n43_w71, 
            w72=> c1_n43_w72, 
            w73=> c1_n43_w73, 
            w74=> c1_n43_w74, 
            w75=> c1_n43_w75, 
            w76=> c1_n43_w76, 
            w77=> c1_n43_w77, 
            w78=> c1_n43_w78, 
            w79=> c1_n43_w79, 
            w80=> c1_n43_w80, 
            w81=> c1_n43_w81, 
            w82=> c1_n43_w82, 
            w83=> c1_n43_w83, 
            w84=> c1_n43_w84, 
            w85=> c1_n43_w85, 
            w86=> c1_n43_w86, 
            w87=> c1_n43_w87, 
            w88=> c1_n43_w88, 
            w89=> c1_n43_w89, 
            w90=> c1_n43_w90, 
            w91=> c1_n43_w91, 
            w92=> c1_n43_w92, 
            w93=> c1_n43_w93, 
            w94=> c1_n43_w94, 
            w95=> c1_n43_w95, 
            w96=> c1_n43_w96, 
            w97=> c1_n43_w97, 
            w98=> c1_n43_w98, 
            w99=> c1_n43_w99, 
            w100=> c1_n43_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n43_y
   );           
            
neuron_inst_44: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n44_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n44_w1, 
            w2=> c1_n44_w2, 
            w3=> c1_n44_w3, 
            w4=> c1_n44_w4, 
            w5=> c1_n44_w5, 
            w6=> c1_n44_w6, 
            w7=> c1_n44_w7, 
            w8=> c1_n44_w8, 
            w9=> c1_n44_w9, 
            w10=> c1_n44_w10, 
            w11=> c1_n44_w11, 
            w12=> c1_n44_w12, 
            w13=> c1_n44_w13, 
            w14=> c1_n44_w14, 
            w15=> c1_n44_w15, 
            w16=> c1_n44_w16, 
            w17=> c1_n44_w17, 
            w18=> c1_n44_w18, 
            w19=> c1_n44_w19, 
            w20=> c1_n44_w20, 
            w21=> c1_n44_w21, 
            w22=> c1_n44_w22, 
            w23=> c1_n44_w23, 
            w24=> c1_n44_w24, 
            w25=> c1_n44_w25, 
            w26=> c1_n44_w26, 
            w27=> c1_n44_w27, 
            w28=> c1_n44_w28, 
            w29=> c1_n44_w29, 
            w30=> c1_n44_w30, 
            w31=> c1_n44_w31, 
            w32=> c1_n44_w32, 
            w33=> c1_n44_w33, 
            w34=> c1_n44_w34, 
            w35=> c1_n44_w35, 
            w36=> c1_n44_w36, 
            w37=> c1_n44_w37, 
            w38=> c1_n44_w38, 
            w39=> c1_n44_w39, 
            w40=> c1_n44_w40, 
            w41=> c1_n44_w41, 
            w42=> c1_n44_w42, 
            w43=> c1_n44_w43, 
            w44=> c1_n44_w44, 
            w45=> c1_n44_w45, 
            w46=> c1_n44_w46, 
            w47=> c1_n44_w47, 
            w48=> c1_n44_w48, 
            w49=> c1_n44_w49, 
            w50=> c1_n44_w50, 
            w51=> c1_n44_w51, 
            w52=> c1_n44_w52, 
            w53=> c1_n44_w53, 
            w54=> c1_n44_w54, 
            w55=> c1_n44_w55, 
            w56=> c1_n44_w56, 
            w57=> c1_n44_w57, 
            w58=> c1_n44_w58, 
            w59=> c1_n44_w59, 
            w60=> c1_n44_w60, 
            w61=> c1_n44_w61, 
            w62=> c1_n44_w62, 
            w63=> c1_n44_w63, 
            w64=> c1_n44_w64, 
            w65=> c1_n44_w65, 
            w66=> c1_n44_w66, 
            w67=> c1_n44_w67, 
            w68=> c1_n44_w68, 
            w69=> c1_n44_w69, 
            w70=> c1_n44_w70, 
            w71=> c1_n44_w71, 
            w72=> c1_n44_w72, 
            w73=> c1_n44_w73, 
            w74=> c1_n44_w74, 
            w75=> c1_n44_w75, 
            w76=> c1_n44_w76, 
            w77=> c1_n44_w77, 
            w78=> c1_n44_w78, 
            w79=> c1_n44_w79, 
            w80=> c1_n44_w80, 
            w81=> c1_n44_w81, 
            w82=> c1_n44_w82, 
            w83=> c1_n44_w83, 
            w84=> c1_n44_w84, 
            w85=> c1_n44_w85, 
            w86=> c1_n44_w86, 
            w87=> c1_n44_w87, 
            w88=> c1_n44_w88, 
            w89=> c1_n44_w89, 
            w90=> c1_n44_w90, 
            w91=> c1_n44_w91, 
            w92=> c1_n44_w92, 
            w93=> c1_n44_w93, 
            w94=> c1_n44_w94, 
            w95=> c1_n44_w95, 
            w96=> c1_n44_w96, 
            w97=> c1_n44_w97, 
            w98=> c1_n44_w98, 
            w99=> c1_n44_w99, 
            w100=> c1_n44_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n44_y
   );           
            
neuron_inst_45: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n45_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n45_w1, 
            w2=> c1_n45_w2, 
            w3=> c1_n45_w3, 
            w4=> c1_n45_w4, 
            w5=> c1_n45_w5, 
            w6=> c1_n45_w6, 
            w7=> c1_n45_w7, 
            w8=> c1_n45_w8, 
            w9=> c1_n45_w9, 
            w10=> c1_n45_w10, 
            w11=> c1_n45_w11, 
            w12=> c1_n45_w12, 
            w13=> c1_n45_w13, 
            w14=> c1_n45_w14, 
            w15=> c1_n45_w15, 
            w16=> c1_n45_w16, 
            w17=> c1_n45_w17, 
            w18=> c1_n45_w18, 
            w19=> c1_n45_w19, 
            w20=> c1_n45_w20, 
            w21=> c1_n45_w21, 
            w22=> c1_n45_w22, 
            w23=> c1_n45_w23, 
            w24=> c1_n45_w24, 
            w25=> c1_n45_w25, 
            w26=> c1_n45_w26, 
            w27=> c1_n45_w27, 
            w28=> c1_n45_w28, 
            w29=> c1_n45_w29, 
            w30=> c1_n45_w30, 
            w31=> c1_n45_w31, 
            w32=> c1_n45_w32, 
            w33=> c1_n45_w33, 
            w34=> c1_n45_w34, 
            w35=> c1_n45_w35, 
            w36=> c1_n45_w36, 
            w37=> c1_n45_w37, 
            w38=> c1_n45_w38, 
            w39=> c1_n45_w39, 
            w40=> c1_n45_w40, 
            w41=> c1_n45_w41, 
            w42=> c1_n45_w42, 
            w43=> c1_n45_w43, 
            w44=> c1_n45_w44, 
            w45=> c1_n45_w45, 
            w46=> c1_n45_w46, 
            w47=> c1_n45_w47, 
            w48=> c1_n45_w48, 
            w49=> c1_n45_w49, 
            w50=> c1_n45_w50, 
            w51=> c1_n45_w51, 
            w52=> c1_n45_w52, 
            w53=> c1_n45_w53, 
            w54=> c1_n45_w54, 
            w55=> c1_n45_w55, 
            w56=> c1_n45_w56, 
            w57=> c1_n45_w57, 
            w58=> c1_n45_w58, 
            w59=> c1_n45_w59, 
            w60=> c1_n45_w60, 
            w61=> c1_n45_w61, 
            w62=> c1_n45_w62, 
            w63=> c1_n45_w63, 
            w64=> c1_n45_w64, 
            w65=> c1_n45_w65, 
            w66=> c1_n45_w66, 
            w67=> c1_n45_w67, 
            w68=> c1_n45_w68, 
            w69=> c1_n45_w69, 
            w70=> c1_n45_w70, 
            w71=> c1_n45_w71, 
            w72=> c1_n45_w72, 
            w73=> c1_n45_w73, 
            w74=> c1_n45_w74, 
            w75=> c1_n45_w75, 
            w76=> c1_n45_w76, 
            w77=> c1_n45_w77, 
            w78=> c1_n45_w78, 
            w79=> c1_n45_w79, 
            w80=> c1_n45_w80, 
            w81=> c1_n45_w81, 
            w82=> c1_n45_w82, 
            w83=> c1_n45_w83, 
            w84=> c1_n45_w84, 
            w85=> c1_n45_w85, 
            w86=> c1_n45_w86, 
            w87=> c1_n45_w87, 
            w88=> c1_n45_w88, 
            w89=> c1_n45_w89, 
            w90=> c1_n45_w90, 
            w91=> c1_n45_w91, 
            w92=> c1_n45_w92, 
            w93=> c1_n45_w93, 
            w94=> c1_n45_w94, 
            w95=> c1_n45_w95, 
            w96=> c1_n45_w96, 
            w97=> c1_n45_w97, 
            w98=> c1_n45_w98, 
            w99=> c1_n45_w99, 
            w100=> c1_n45_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n45_y
   );           
            
neuron_inst_46: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n46_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n46_w1, 
            w2=> c1_n46_w2, 
            w3=> c1_n46_w3, 
            w4=> c1_n46_w4, 
            w5=> c1_n46_w5, 
            w6=> c1_n46_w6, 
            w7=> c1_n46_w7, 
            w8=> c1_n46_w8, 
            w9=> c1_n46_w9, 
            w10=> c1_n46_w10, 
            w11=> c1_n46_w11, 
            w12=> c1_n46_w12, 
            w13=> c1_n46_w13, 
            w14=> c1_n46_w14, 
            w15=> c1_n46_w15, 
            w16=> c1_n46_w16, 
            w17=> c1_n46_w17, 
            w18=> c1_n46_w18, 
            w19=> c1_n46_w19, 
            w20=> c1_n46_w20, 
            w21=> c1_n46_w21, 
            w22=> c1_n46_w22, 
            w23=> c1_n46_w23, 
            w24=> c1_n46_w24, 
            w25=> c1_n46_w25, 
            w26=> c1_n46_w26, 
            w27=> c1_n46_w27, 
            w28=> c1_n46_w28, 
            w29=> c1_n46_w29, 
            w30=> c1_n46_w30, 
            w31=> c1_n46_w31, 
            w32=> c1_n46_w32, 
            w33=> c1_n46_w33, 
            w34=> c1_n46_w34, 
            w35=> c1_n46_w35, 
            w36=> c1_n46_w36, 
            w37=> c1_n46_w37, 
            w38=> c1_n46_w38, 
            w39=> c1_n46_w39, 
            w40=> c1_n46_w40, 
            w41=> c1_n46_w41, 
            w42=> c1_n46_w42, 
            w43=> c1_n46_w43, 
            w44=> c1_n46_w44, 
            w45=> c1_n46_w45, 
            w46=> c1_n46_w46, 
            w47=> c1_n46_w47, 
            w48=> c1_n46_w48, 
            w49=> c1_n46_w49, 
            w50=> c1_n46_w50, 
            w51=> c1_n46_w51, 
            w52=> c1_n46_w52, 
            w53=> c1_n46_w53, 
            w54=> c1_n46_w54, 
            w55=> c1_n46_w55, 
            w56=> c1_n46_w56, 
            w57=> c1_n46_w57, 
            w58=> c1_n46_w58, 
            w59=> c1_n46_w59, 
            w60=> c1_n46_w60, 
            w61=> c1_n46_w61, 
            w62=> c1_n46_w62, 
            w63=> c1_n46_w63, 
            w64=> c1_n46_w64, 
            w65=> c1_n46_w65, 
            w66=> c1_n46_w66, 
            w67=> c1_n46_w67, 
            w68=> c1_n46_w68, 
            w69=> c1_n46_w69, 
            w70=> c1_n46_w70, 
            w71=> c1_n46_w71, 
            w72=> c1_n46_w72, 
            w73=> c1_n46_w73, 
            w74=> c1_n46_w74, 
            w75=> c1_n46_w75, 
            w76=> c1_n46_w76, 
            w77=> c1_n46_w77, 
            w78=> c1_n46_w78, 
            w79=> c1_n46_w79, 
            w80=> c1_n46_w80, 
            w81=> c1_n46_w81, 
            w82=> c1_n46_w82, 
            w83=> c1_n46_w83, 
            w84=> c1_n46_w84, 
            w85=> c1_n46_w85, 
            w86=> c1_n46_w86, 
            w87=> c1_n46_w87, 
            w88=> c1_n46_w88, 
            w89=> c1_n46_w89, 
            w90=> c1_n46_w90, 
            w91=> c1_n46_w91, 
            w92=> c1_n46_w92, 
            w93=> c1_n46_w93, 
            w94=> c1_n46_w94, 
            w95=> c1_n46_w95, 
            w96=> c1_n46_w96, 
            w97=> c1_n46_w97, 
            w98=> c1_n46_w98, 
            w99=> c1_n46_w99, 
            w100=> c1_n46_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n46_y
   );           
            
neuron_inst_47: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n47_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n47_w1, 
            w2=> c1_n47_w2, 
            w3=> c1_n47_w3, 
            w4=> c1_n47_w4, 
            w5=> c1_n47_w5, 
            w6=> c1_n47_w6, 
            w7=> c1_n47_w7, 
            w8=> c1_n47_w8, 
            w9=> c1_n47_w9, 
            w10=> c1_n47_w10, 
            w11=> c1_n47_w11, 
            w12=> c1_n47_w12, 
            w13=> c1_n47_w13, 
            w14=> c1_n47_w14, 
            w15=> c1_n47_w15, 
            w16=> c1_n47_w16, 
            w17=> c1_n47_w17, 
            w18=> c1_n47_w18, 
            w19=> c1_n47_w19, 
            w20=> c1_n47_w20, 
            w21=> c1_n47_w21, 
            w22=> c1_n47_w22, 
            w23=> c1_n47_w23, 
            w24=> c1_n47_w24, 
            w25=> c1_n47_w25, 
            w26=> c1_n47_w26, 
            w27=> c1_n47_w27, 
            w28=> c1_n47_w28, 
            w29=> c1_n47_w29, 
            w30=> c1_n47_w30, 
            w31=> c1_n47_w31, 
            w32=> c1_n47_w32, 
            w33=> c1_n47_w33, 
            w34=> c1_n47_w34, 
            w35=> c1_n47_w35, 
            w36=> c1_n47_w36, 
            w37=> c1_n47_w37, 
            w38=> c1_n47_w38, 
            w39=> c1_n47_w39, 
            w40=> c1_n47_w40, 
            w41=> c1_n47_w41, 
            w42=> c1_n47_w42, 
            w43=> c1_n47_w43, 
            w44=> c1_n47_w44, 
            w45=> c1_n47_w45, 
            w46=> c1_n47_w46, 
            w47=> c1_n47_w47, 
            w48=> c1_n47_w48, 
            w49=> c1_n47_w49, 
            w50=> c1_n47_w50, 
            w51=> c1_n47_w51, 
            w52=> c1_n47_w52, 
            w53=> c1_n47_w53, 
            w54=> c1_n47_w54, 
            w55=> c1_n47_w55, 
            w56=> c1_n47_w56, 
            w57=> c1_n47_w57, 
            w58=> c1_n47_w58, 
            w59=> c1_n47_w59, 
            w60=> c1_n47_w60, 
            w61=> c1_n47_w61, 
            w62=> c1_n47_w62, 
            w63=> c1_n47_w63, 
            w64=> c1_n47_w64, 
            w65=> c1_n47_w65, 
            w66=> c1_n47_w66, 
            w67=> c1_n47_w67, 
            w68=> c1_n47_w68, 
            w69=> c1_n47_w69, 
            w70=> c1_n47_w70, 
            w71=> c1_n47_w71, 
            w72=> c1_n47_w72, 
            w73=> c1_n47_w73, 
            w74=> c1_n47_w74, 
            w75=> c1_n47_w75, 
            w76=> c1_n47_w76, 
            w77=> c1_n47_w77, 
            w78=> c1_n47_w78, 
            w79=> c1_n47_w79, 
            w80=> c1_n47_w80, 
            w81=> c1_n47_w81, 
            w82=> c1_n47_w82, 
            w83=> c1_n47_w83, 
            w84=> c1_n47_w84, 
            w85=> c1_n47_w85, 
            w86=> c1_n47_w86, 
            w87=> c1_n47_w87, 
            w88=> c1_n47_w88, 
            w89=> c1_n47_w89, 
            w90=> c1_n47_w90, 
            w91=> c1_n47_w91, 
            w92=> c1_n47_w92, 
            w93=> c1_n47_w93, 
            w94=> c1_n47_w94, 
            w95=> c1_n47_w95, 
            w96=> c1_n47_w96, 
            w97=> c1_n47_w97, 
            w98=> c1_n47_w98, 
            w99=> c1_n47_w99, 
            w100=> c1_n47_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n47_y
   );           
            
neuron_inst_48: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n48_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n48_w1, 
            w2=> c1_n48_w2, 
            w3=> c1_n48_w3, 
            w4=> c1_n48_w4, 
            w5=> c1_n48_w5, 
            w6=> c1_n48_w6, 
            w7=> c1_n48_w7, 
            w8=> c1_n48_w8, 
            w9=> c1_n48_w9, 
            w10=> c1_n48_w10, 
            w11=> c1_n48_w11, 
            w12=> c1_n48_w12, 
            w13=> c1_n48_w13, 
            w14=> c1_n48_w14, 
            w15=> c1_n48_w15, 
            w16=> c1_n48_w16, 
            w17=> c1_n48_w17, 
            w18=> c1_n48_w18, 
            w19=> c1_n48_w19, 
            w20=> c1_n48_w20, 
            w21=> c1_n48_w21, 
            w22=> c1_n48_w22, 
            w23=> c1_n48_w23, 
            w24=> c1_n48_w24, 
            w25=> c1_n48_w25, 
            w26=> c1_n48_w26, 
            w27=> c1_n48_w27, 
            w28=> c1_n48_w28, 
            w29=> c1_n48_w29, 
            w30=> c1_n48_w30, 
            w31=> c1_n48_w31, 
            w32=> c1_n48_w32, 
            w33=> c1_n48_w33, 
            w34=> c1_n48_w34, 
            w35=> c1_n48_w35, 
            w36=> c1_n48_w36, 
            w37=> c1_n48_w37, 
            w38=> c1_n48_w38, 
            w39=> c1_n48_w39, 
            w40=> c1_n48_w40, 
            w41=> c1_n48_w41, 
            w42=> c1_n48_w42, 
            w43=> c1_n48_w43, 
            w44=> c1_n48_w44, 
            w45=> c1_n48_w45, 
            w46=> c1_n48_w46, 
            w47=> c1_n48_w47, 
            w48=> c1_n48_w48, 
            w49=> c1_n48_w49, 
            w50=> c1_n48_w50, 
            w51=> c1_n48_w51, 
            w52=> c1_n48_w52, 
            w53=> c1_n48_w53, 
            w54=> c1_n48_w54, 
            w55=> c1_n48_w55, 
            w56=> c1_n48_w56, 
            w57=> c1_n48_w57, 
            w58=> c1_n48_w58, 
            w59=> c1_n48_w59, 
            w60=> c1_n48_w60, 
            w61=> c1_n48_w61, 
            w62=> c1_n48_w62, 
            w63=> c1_n48_w63, 
            w64=> c1_n48_w64, 
            w65=> c1_n48_w65, 
            w66=> c1_n48_w66, 
            w67=> c1_n48_w67, 
            w68=> c1_n48_w68, 
            w69=> c1_n48_w69, 
            w70=> c1_n48_w70, 
            w71=> c1_n48_w71, 
            w72=> c1_n48_w72, 
            w73=> c1_n48_w73, 
            w74=> c1_n48_w74, 
            w75=> c1_n48_w75, 
            w76=> c1_n48_w76, 
            w77=> c1_n48_w77, 
            w78=> c1_n48_w78, 
            w79=> c1_n48_w79, 
            w80=> c1_n48_w80, 
            w81=> c1_n48_w81, 
            w82=> c1_n48_w82, 
            w83=> c1_n48_w83, 
            w84=> c1_n48_w84, 
            w85=> c1_n48_w85, 
            w86=> c1_n48_w86, 
            w87=> c1_n48_w87, 
            w88=> c1_n48_w88, 
            w89=> c1_n48_w89, 
            w90=> c1_n48_w90, 
            w91=> c1_n48_w91, 
            w92=> c1_n48_w92, 
            w93=> c1_n48_w93, 
            w94=> c1_n48_w94, 
            w95=> c1_n48_w95, 
            w96=> c1_n48_w96, 
            w97=> c1_n48_w97, 
            w98=> c1_n48_w98, 
            w99=> c1_n48_w99, 
            w100=> c1_n48_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n48_y
   );           
            
neuron_inst_49: ENTITY work.neuron_comb_ReLU_100n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n49_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n49_w1, 
            w2=> c1_n49_w2, 
            w3=> c1_n49_w3, 
            w4=> c1_n49_w4, 
            w5=> c1_n49_w5, 
            w6=> c1_n49_w6, 
            w7=> c1_n49_w7, 
            w8=> c1_n49_w8, 
            w9=> c1_n49_w9, 
            w10=> c1_n49_w10, 
            w11=> c1_n49_w11, 
            w12=> c1_n49_w12, 
            w13=> c1_n49_w13, 
            w14=> c1_n49_w14, 
            w15=> c1_n49_w15, 
            w16=> c1_n49_w16, 
            w17=> c1_n49_w17, 
            w18=> c1_n49_w18, 
            w19=> c1_n49_w19, 
            w20=> c1_n49_w20, 
            w21=> c1_n49_w21, 
            w22=> c1_n49_w22, 
            w23=> c1_n49_w23, 
            w24=> c1_n49_w24, 
            w25=> c1_n49_w25, 
            w26=> c1_n49_w26, 
            w27=> c1_n49_w27, 
            w28=> c1_n49_w28, 
            w29=> c1_n49_w29, 
            w30=> c1_n49_w30, 
            w31=> c1_n49_w31, 
            w32=> c1_n49_w32, 
            w33=> c1_n49_w33, 
            w34=> c1_n49_w34, 
            w35=> c1_n49_w35, 
            w36=> c1_n49_w36, 
            w37=> c1_n49_w37, 
            w38=> c1_n49_w38, 
            w39=> c1_n49_w39, 
            w40=> c1_n49_w40, 
            w41=> c1_n49_w41, 
            w42=> c1_n49_w42, 
            w43=> c1_n49_w43, 
            w44=> c1_n49_w44, 
            w45=> c1_n49_w45, 
            w46=> c1_n49_w46, 
            w47=> c1_n49_w47, 
            w48=> c1_n49_w48, 
            w49=> c1_n49_w49, 
            w50=> c1_n49_w50, 
            w51=> c1_n49_w51, 
            w52=> c1_n49_w52, 
            w53=> c1_n49_w53, 
            w54=> c1_n49_w54, 
            w55=> c1_n49_w55, 
            w56=> c1_n49_w56, 
            w57=> c1_n49_w57, 
            w58=> c1_n49_w58, 
            w59=> c1_n49_w59, 
            w60=> c1_n49_w60, 
            w61=> c1_n49_w61, 
            w62=> c1_n49_w62, 
            w63=> c1_n49_w63, 
            w64=> c1_n49_w64, 
            w65=> c1_n49_w65, 
            w66=> c1_n49_w66, 
            w67=> c1_n49_w67, 
            w68=> c1_n49_w68, 
            w69=> c1_n49_w69, 
            w70=> c1_n49_w70, 
            w71=> c1_n49_w71, 
            w72=> c1_n49_w72, 
            w73=> c1_n49_w73, 
            w74=> c1_n49_w74, 
            w75=> c1_n49_w75, 
            w76=> c1_n49_w76, 
            w77=> c1_n49_w77, 
            w78=> c1_n49_w78, 
            w79=> c1_n49_w79, 
            w80=> c1_n49_w80, 
            w81=> c1_n49_w81, 
            w82=> c1_n49_w82, 
            w83=> c1_n49_w83, 
            w84=> c1_n49_w84, 
            w85=> c1_n49_w85, 
            w86=> c1_n49_w86, 
            w87=> c1_n49_w87, 
            w88=> c1_n49_w88, 
            w89=> c1_n49_w89, 
            w90=> c1_n49_w90, 
            w91=> c1_n49_w91, 
            w92=> c1_n49_w92, 
            w93=> c1_n49_w93, 
            w94=> c1_n49_w94, 
            w95=> c1_n49_w95, 
            w96=> c1_n49_w96, 
            w97=> c1_n49_w97, 
            w98=> c1_n49_w98, 
            w99=> c1_n49_w99, 
            w100=> c1_n49_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n49_y
   );           
             
END ARCHITECTURE;
