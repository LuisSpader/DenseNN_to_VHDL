
--https://stackoverflow.com/questions/17579716/implementing-rom-in-xilinx-vhdl
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
----------------
ENTITY ROM_Sigmoid_8bit IS
	GENERIC (
		addr_width : INTEGER := 256; -- store 256 elements
		addr_bits  : INTEGER := 8;   -- required bits to store 256 elements
		data_width : INTEGER := 8    -- each element has 8-bits
	);
	PORT (
		address  : IN STD_LOGIC_VECTOR(addr_bits - 1 DOWNTO 0);
		data_out : OUT STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0)
	);
END ENTITY;
------------------
ARCHITECTURE arch OF ROM_Sigmoid_8bit IS
	TYPE memory IS ARRAY (0 TO addr_width - 1) OF STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0);
	CONSTANT myrom : memory := (
		--"int_f_x",--(address)  =integer_MAC|| f(x)               = int_f_x 
		"10000000", -- (00000000) = 0.0       || 128.0              = 128.0
		"10000010", -- (00000001) = 1.0       || 130.79955347088494 = 130.0
		"10000101", -- (00000010) = 2.0       || 133.59642981673    = 133.0
		"10001000", -- (00000011) = 3.0       || 136.38796214291455 = 136.0
		"10001011", -- (00000100) = 4.0       || 139.1715039326922  = 139.0
		"10001101", -- (00000101) = 5.0       || 141.9444390298694  = 141.0
		"10010000", -- (00000110) = 6.0       || 144.70419137717758 = 144.0
		"10010011", -- (00000111) = 7.0       || 147.44823443416874 = 147.0
		"10010110", -- (00001000) = 8.0       || 150.1741002028365  = 150.0
		"10011000", -- (00001001) = 9.0       || 152.8793877944536  = 152.0
		"10011011", -- (00001010) = 10.0      || 155.56177147722028 = 155.0
		"10011110", -- (00001011) = 11.0      || 158.21900815110592 = 158.0
		"10100000", -- (00001100) = 12.0      || 160.84894420361377 = 160.0
		"10100011", -- (00001101) = 13.0      || 163.4495217079567  = 163.0
		"10100110", -- (00001110) = 14.0      || 166.01878393316375 = 166.0
		"10101000", -- (00001111) = 15.0      || 168.55488014379085 = 168.0
		"10101011", -- (00010000) = 16.0      || 171.05606967505054 = 171.0
		"10101101", -- (00010001) = 17.0      || 173.52072527716751 = 173.0
		"10101111", -- (00010010) = 18.0      || 175.94733573048427 = 175.0
		"10110010", -- (00010011) = 19.0      || 178.3345077401747  = 178.0
		"10110100", -- (00010100) = 20.0      || 180.68096712627488 = 180.0
		"10110110", -- (00010101) = 21.0      || 182.98555933102264 = 182.0
		"10111001", -- (00010110) = 22.0      || 185.24724927115267 = 185.0
		"10111011", -- (00010111) = 23.0      || 187.46512056776362 = 187.0
		"10111101", -- (00011000) = 24.0      || 189.6383741906314  = 189.0
		"10111111", -- (00011001) = 25.0      || 191.76632655737023 = 191.0
		"11000001", -- (00011010) = 26.0      || 193.84840713063423 = 193.0
		"11000011", -- (00011011) = 27.0      || 195.88415555862744 = 195.0
		"11000101", -- (00011100) = 28.0      || 197.87321840556507 = 197.0
		"11000111", -- (00011101) = 29.0      || 199.8153455194442  = 199.0
		"11001001", -- (00011110) = 30.0      || 201.71038608458105 = 201.0
		"11001011", -- (00011111) = 31.0      || 203.55828440590156 = 203.0
		"11001101", -- (00100000) = 32.0      || 205.3590754709969  = 205.0
		"11001111", -- (00100001) = 33.0      || 207.1128803345236  = 207.0
		"11010000", -- (00100010) = 34.0      || 208.819901367714   = 208.0
		"11010010", -- (00100011) = 35.0      || 210.48041741361928 = 210.0
		"11010100", -- (00100100) = 36.0      || 212.09477888629738 = 212.0
		"11010101", -- (00100101) = 37.0      || 213.66340284954757 = 213.0
		"11010111", -- (00100110) = 38.0      || 215.1867681080277  = 215.0
		"11011000", -- (00100111) = 39.0      || 216.66541034073072 = 216.0
		"11011010", -- (00101000) = 40.0      || 218.0999173038875  = 218.0
		"11011011", -- (00101001) = 41.0      || 219.49092412744895 = 219.0
		"11011100", -- (00101010) = 42.0      || 220.8391087264176  = 220.0
		"11011110", -- (00101011) = 43.0      || 222.1451873454842  = 222.0
		"11011111", -- (00101100) = 44.0      || 223.40991025270483 = 223.0
		"11100000", -- (00101101) = 45.0      || 224.6340575953512  = 224.0
		"11100001", -- (00101110) = 46.0      || 225.8184354286031  = 225.0
		"11100010", -- (00101111) = 47.0      || 226.96387192543793 = 226.0
		"11100100", -- (00110000) = 48.0      || 228.0712137739231  = 228.0
		"11100101", -- (00110001) = 49.0      || 229.14132276613313 = 229.0
		"11100110", -- (00110010) = 50.0      || 230.17507258110555 = 230.0
		"11100111", -- (00110011) = 51.0      || 231.17334576261152 = 231.0
		"11101000", -- (00110100) = 52.0      || 232.13703089105314 = 232.0
		"11101001", -- (00110101) = 53.0      || 233.0670199474983  = 233.0
		"11101001", -- (00110110) = 54.0      || 233.9642058667285  = 233.0
		"11101010", -- (00110111) = 55.0      || 234.82948027519006 = 234.0
		"11101011", -- (00111000) = 56.0      || 235.66373140890153 = 235.0
		"11101100", -- (00111001) = 57.0      || 236.4678422056685  = 236.0
		"11101101", -- (00111010) = 58.0      || 237.24268856538296 = 237.0
		"11101101", -- (00111011) = 59.0      || 237.9891377717278  = 237.0
		"11101110", -- (00111100) = 60.0      || 238.70804706825496 = 238.0
		"11101111", -- (00111101) = 61.0      || 239.40026238155605 = 239.0
		"11110000", -- (00111110) = 62.0      || 240.06661718407545 = 240.0
		"11110000", -- (00111111) = 63.0      || 240.7079314890315  = 240.0
		"11110001", -- (01000000) = 64.0      || 241.3250109698896  = 241.0
		"11110001", -- (01000001) = 65.0      || 241.91864619687576 = 241.0
		"11110010", -- (01000010) = 66.0      || 242.48961198310965 = 242.0
		"11110011", -- (01000011) = 67.0      || 243.03866683307706 = 243.0
		"11110011", -- (01000100) = 68.0      || 243.56655248633442 = 243.0
		"11110100", -- (01000101) = 69.0      || 244.07399354954848 = 244.0
		"11110100", -- (01000110) = 70.0      || 244.56169721020154 = 244.0
		"11110101", -- (01000111) = 71.0      || 245.03035302554926 = 245.0
		"11110101", -- (01001000) = 72.0      || 245.48063278068096 = 245.0
		"11110101", -- (01001001) = 73.0      || 245.9131904098127  = 245.0
		"11110110", -- (01001010) = 74.0      || 246.3286619752277  = 246.0
		"11110110", -- (01001011) = 75.0      || 246.72766569856648 = 246.0
		"11110111", -- (01001100) = 76.0      || 247.11080203946045 = 247.0
		"11110111", -- (01001101) = 77.0      || 247.47865381678946 = 247.0
		"11110111", -- (01001110) = 78.0      || 247.8317863681286  = 247.0
		"11111000", -- (01001111) = 79.0      || 248.17074774322967 = 248.0
		"11111000", -- (01010000) = 80.0      || 248.49606892765277 = 248.0
		"11111000", -- (01010001) = 81.0      || 248.80826409293064 = 248.0
		"11111001", -- (01010010) = 82.0      || 249.10783086989977 = 249.0
		"11111001", -- (01010011) = 83.0      || 249.3952506420807  = 249.0
		"11111001", -- (01010100) = 84.0      || 249.67098885622383 = 249.0
		"11111001", -- (01010101) = 85.0      || 249.93549534736016 = 249.0
		"11111010", -- (01010110) = 86.0      || 250.18920467591147 = 250.0
		"11111010", -- (01010111) = 87.0      || 250.4325364746162  = 250.0
		"11111010", -- (01011000) = 88.0      || 250.6658958032178  = 250.0
		"11111010", -- (01011001) = 89.0      || 250.88967350904375 = 250.0
		"11111011", -- (01011010) = 90.0      || 251.10424659177247 = 251.0
		"11111011", -- (01011011) = 91.0      || 251.30997857084472 = 251.0
		"11111011", -- (01011100) = 92.0      || 251.50721985412497 = 251.0
		"11111011", -- (01011101) = 93.0      || 251.6963081065567  = 251.0
		"11111011", -- (01011110) = 94.0      || 251.87756861768625 = 251.0
		"11111100", -- (01011111) = 95.0      || 252.05131466704864 = 252.0
		"11111100", -- (01100000) = 96.0      || 252.2178478865221  = 252.0
		"11111100", -- (01100001) = 97.0      || 252.3774586188595  = 252.0
		"11111100", -- (01100010) = 98.0      || 252.53042627170205 = 252.0
		"11111100", -- (01100011) = 99.0      || 252.6770196664673  = 252.0
		"11111100", -- (01100100) = 100.0     || 252.81749738158442 = 252.0
		"11111100", -- (01100101) = 101.0     || 252.95210808962463 = 252.0
		"11111101", -- (01100110) = 102.0     || 253.08109088794197 = 253.0
		"11111101", -- (01100111) = 103.0     || 253.20467562250147 = 253.0
		"11111101", -- (01101000) = 104.0     || 253.32308320462894 = 253.0
		"11111101", -- (01101001) = 105.0     || 253.43652592046766 = 253.0
		"11111101", -- (01101010) = 106.0     || 253.54520773297327 = 253.0
		"11111101", -- (01101011) = 107.0     || 253.64932457632193 = 253.0
		"11111101", -- (01101100) = 108.0     || 253.74906464264322 = 253.0
		"11111101", -- (01101101) = 109.0     || 253.84460866102432 = 253.0
		"11111101", -- (01101110) = 110.0     || 253.93613016876247 = 253.0
		"11111110", -- (01101111) = 111.0     || 254.0237957748705  = 254.0
		"11111110", -- (01110000) = 112.0     || 254.10776541586384 = 254.0
		"11111110", -- (01110001) = 113.0     || 254.18819260387994 = 254.0
		"11111110", -- (01110010) = 114.0     || 254.26522466719953 = 254.0
		"11111110", -- (01110011) = 115.0     || 254.3390029832559  = 254.0
		"11111110", -- (01110100) = 116.0     || 254.40966320423354 = 254.0
		"11111110", -- (01110101) = 117.0     || 254.47733547536947 = 254.0
		"11111110", -- (01110110) = 118.0     || 254.54214464608148 = 254.0
		"11111110", -- (01110111) = 119.0     || 254.60421047405794 = 254.0
		"11111110", -- (01111000) = 120.0     || 254.66364782244906 = 254.0
		"11111110", -- (01111001) = 121.0     || 254.72056685030938 = 254.0
		"11111110", -- (01111010) = 122.0     || 254.775073196443   = 254.0
		"11111110", -- (01111011) = 123.0     || 254.82726815680954 = 254.0
		"11111110", -- (01111100) = 124.0     || 254.87724885565115 = 254.0
		"11111110", -- (01111101) = 125.0     || 254.92510841050319 = 254.0
		"11111110", -- (01111110) = 126.0     || 254.97093609125218 = 254.0
		"11111111", -- (01111111) = 127.0     || 255.01481747340657 = 255.0
		"00000000", -- (10000000) = -128.0    || 0.9431654142556132 = 0.0
		"00000000", -- (10000001) = -127.0    || 0.9851825265934124 = 0.0
		"00000001", -- (10000010) = -126.0    || 1.0290639087477775 = 1.0
		"00000001", -- (10000011) = -125.0    || 1.0748915894967983 = 1.0
		"00000001", -- (10000100) = -124.0    || 1.1227511443488492 = 1.0
		"00000001", -- (10000101) = -123.0    || 1.1727318431904823 = 1.0
		"00000001", -- (10000110) = -122.0    || 1.2249268035570005 = 1.0
		"00000001", -- (10000111) = -121.0    || 1.2794331496906086 = 1.0
		"00000001", -- (10001000) = -120.0    || 1.3363521775509497 = 1.0
		"00000001", -- (10001001) = -119.0    || 1.3957895259420845 = 1.0
		"00000001", -- (10001010) = -118.0    || 1.457855353918504  = 1.0
		"00000001", -- (10001011) = -117.0    || 1.5226645246305492 = 1.0
		"00000001", -- (10001100) = -116.0    || 1.590336795766455  = 1.0
		"00000001", -- (10001101) = -115.0    || 1.6609970167441164 = 1.0
		"00000001", -- (10001110) = -114.0    || 1.73477533280049   = 1.0
		"00000001", -- (10001111) = -113.0    || 1.811807396120073  = 1.0
		"00000001", -- (10010000) = -112.0    || 1.892234584136186  = 1.0
		"00000001", -- (10010001) = -111.0    || 1.9762042251295215 = 1.0
		"00000010", -- (10010010) = -110.0    || 2.06386983123754   = 2.0
		"00000010", -- (10010011) = -109.0    || 2.155391338975693  = 2.0
		"00000010", -- (10010100) = -108.0    || 2.2509353573567803 = 2.0
		"00000010", -- (10010101) = -107.0    || 2.3506754236780787 = 2.0
		"00000010", -- (10010110) = -106.0    || 2.454792267026737  = 2.0
		"00000010", -- (10010111) = -105.0    || 2.563474079532323  = 2.0
		"00000010", -- (10011000) = -104.0    || 2.6769167953710262 = 2.0
		"00000010", -- (10011001) = -103.0    || 2.7953243774985372 = 2.0
		"00000010", -- (10011010) = -102.0    || 2.9189091120580306 = 2.0
		"00000011", -- (10011011) = -101.0    || 3.0478919103753572 = 3.0
		"00000011", -- (10011100) = -100.0    || 3.18250261841557   = 3.0
		"00000011", -- (10011101) = -99.0     || 3.3229803335326857 = 3.0
		"00000011", -- (10011110) = -98.0     || 3.4695737282979517 = 3.0
		"00000011", -- (10011111) = -97.0     || 3.6225413811405303 = 3.0
		"00000011", -- (10100000) = -96.0     || 3.7821521134779053 = 3.0
		"00000011", -- (10100001) = -95.0     || 3.948685332951331  = 3.0
		"00000100", -- (10100010) = -94.0     || 4.122431382313737  = 4.0
		"00000100", -- (10100011) = -93.0     || 4.303691893443283  = 4.0
		"00000100", -- (10100100) = -92.0     || 4.492780145875043  = 4.0
		"00000100", -- (10100101) = -91.0     || 4.690021429155295  = 4.0
		"00000100", -- (10100110) = -90.0     || 4.895753408227562  = 4.0
		"00000101", -- (10100111) = -89.0     || 5.110326490956257  = 5.0
		"00000101", -- (10101000) = -88.0     || 5.3341041967821905 = 5.0
		"00000101", -- (10101001) = -87.0     || 5.567463525383797  = 5.0
		"00000101", -- (10101010) = -86.0     || 5.81079532408854   = 5.0
		"00000110", -- (10101011) = -85.0     || 6.064504652639856  = 6.0
		"00000110", -- (10101100) = -84.0     || 6.3290111437761585 = 6.0
		"00000110", -- (10101101) = -83.0     || 6.604749357919308  = 6.0
		"00000110", -- (10101110) = -82.0     || 6.892169130100257  = 6.0
		"00000111", -- (10101111) = -81.0     || 7.191735907069339  = 7.0
		"00000111", -- (10110000) = -80.0     || 7.503931072347218  = 7.0
		"00000111", -- (10110001) = -79.0     || 7.829252256770357  = 7.0
		"00001000", -- (10110010) = -78.0     || 8.168213631871376  = 8.0
		"00001000", -- (10110011) = -77.0     || 8.521346183210536  = 8.0
		"00001000", -- (10110100) = -76.0     || 8.889197960539537  = 8.0
		"00001001", -- (10110101) = -75.0     || 9.272334301433533  = 9.0
		"00001001", -- (10110110) = -74.0     || 9.67133802477231   = 9.0
		"00001010", -- (10110111) = -73.0     || 10.086809590187293 = 10.0
		"00001010", -- (10111000) = -72.0     || 10.519367219319044 = 10.0
		"00001010", -- (10111001) = -71.0     || 10.969646974450724 = 10.0
		"00001011", -- (10111010) = -70.0     || 11.438302789798453 = 11.0
		"00001011", -- (10111011) = -69.0     || 11.926006450451535 = 11.0
		"00001100", -- (10111100) = -68.0     || 12.43344751366557  = 12.0
		"00001100", -- (10111101) = -67.0     || 12.961333166922968 = 12.0
		"00001101", -- (10111110) = -66.0     || 13.510388016890333 = 13.0
		"00001110", -- (10111111) = -65.0     || 14.08135380312426  = 14.0
		"00001110", -- (11000000) = -64.0     || 14.674989030110401 = 14.0
		"00001111", -- (11000001) = -63.0     || 15.292068510968507 = 15.0
		"00001111", -- (11000010) = -62.0     || 15.933382815924531 = 15.0
		"00010000", -- (11000011) = -61.0     || 16.59973761844398  = 16.0
		"00010001", -- (11000100) = -60.0     || 17.29195293174505  = 17.0
		"00010010", -- (11000101) = -59.0     || 18.01086222827223  = 18.0
		"00010010", -- (11000110) = -58.0     || 18.757311434617044 = 18.0
		"00010011", -- (11000111) = -57.0     || 19.532157794331532 = 19.0
		"00010100", -- (11001000) = -56.0     || 20.33626859109847  = 20.0
		"00010101", -- (11001001) = -55.0     || 21.170519724809946 = 21.0
		"00010110", -- (11001010) = -54.0     || 22.035794133271526 = 22.0
		"00010110", -- (11001011) = -53.0     || 22.93298005250171  = 22.0
		"00010111", -- (11001100) = -52.0     || 23.862969108946842 = 23.0
		"00011000", -- (11001101) = -51.0     || 24.826654237388475 = 24.0
		"00011001", -- (11001110) = -50.0     || 25.824927418894468 = 25.0
		"00011010", -- (11001111) = -49.0     || 26.858677233866867 = 26.0
		"00011011", -- (11010000) = -48.0     || 27.928786226076923 = 27.0
		"00011101", -- (11010001) = -47.0     || 29.036128074562075 = 29.0
		"00011110", -- (11010010) = -46.0     || 30.181564571396905 = 30.0
		"00011111", -- (11010011) = -45.0     || 31.36594240464876  = 31.0
		"00100000", -- (11010100) = -44.0     || 32.59008974729516  = 32.0
		"00100001", -- (11010101) = -43.0     || 33.8548126545158   = 33.0
		"00100011", -- (11010110) = -42.0     || 35.1608912735824   = 35.0
		"00100100", -- (11010111) = -41.0     || 36.509075872551044 = 36.0
		"00100101", -- (11011000) = -40.0     || 37.900082696112506 = 37.0
		"00100111", -- (11011001) = -39.0     || 39.33458965926929  = 39.0
		"00101000", -- (11011010) = -38.0     || 40.813231891972286 = 40.0
		"00101010", -- (11011011) = -37.0     || 42.336597150452434 = 42.0
		"00101011", -- (11011100) = -36.0     || 43.90522111370262  = 43.0
		"00101101", -- (11011101) = -35.0     || 45.51958258638069  = 45.0
		"00101111", -- (11011110) = -34.0     || 47.18009863228597  = 47.0
		"00110000", -- (11011111) = -33.0     || 48.88711966547641  = 48.0
		"00110010", -- (11100000) = -32.0     || 50.64092452900307  = 50.0
		"00110100", -- (11100001) = -31.0     || 52.441715594098426 = 52.0
		"00110110", -- (11100010) = -30.0     || 54.28961391541896  = 54.0
		"00111000", -- (11100011) = -29.0     || 56.184654480555785 = 56.0
		"00111010", -- (11100100) = -28.0     || 58.126781594434945 = 58.0
		"00111100", -- (11100101) = -27.0     || 60.11584444137255  = 60.0
		"00111110", -- (11100110) = -26.0     || 62.15159286936576  = 62.0
		"01000000", -- (11100111) = -25.0     || 64.23367344262975  = 64.0
		"01000010", -- (11101000) = -24.0     || 66.36162580936859  = 66.0
		"01000100", -- (11101001) = -23.0     || 68.5348794322364   = 68.0
		"01000110", -- (11101010) = -22.0     || 70.75275072884732  = 70.0
		"01001001", -- (11101011) = -21.0     || 73.01444066897737  = 73.0
		"01001011", -- (11101100) = -20.0     || 75.31903287372512  = 75.0
		"01001101", -- (11101101) = -19.0     || 77.6654922598253   = 77.0
		"01010000", -- (11101110) = -18.0     || 80.05266426951576  = 80.0
		"01010010", -- (11101111) = -17.0     || 82.47927472283249  = 82.0
		"01010100", -- (11110000) = -16.0     || 84.94393032494948  = 84.0
		"01010111", -- (11110001) = -15.0     || 87.44511985620915  = 87.0
		"01011001", -- (11110010) = -14.0     || 89.98121606683623  = 89.0
		"01011100", -- (11110011) = -13.0     || 92.55047829204331  = 92.0
		"01011111", -- (11110100) = -12.0     || 95.15105579638626  = 95.0
		"01100001", -- (11110101) = -11.0     || 97.78099184889408  = 97.0
		"01100100", -- (11110110) = -10.0     || 100.43822852277974 = 100.0
		"01100111", -- (11110111) = -9.0      || 103.12061220554642 = 103.0
		"01101001", -- (11111000) = -8.0      || 105.82589979716352 = 105.0
		"01101100", -- (11111001) = -7.0      || 108.55176556583123 = 108.0
		"01101111", -- (11111010) = -6.0      || 111.29580862282243 = 111.0
		"01110010", -- (11111011) = -5.0      || 114.05556097013061 = 114.0
		"01110100", -- (11111100) = -4.0      || 116.82849606730782 = 116.0
		"01110111", -- (11111101) = -3.0      || 119.61203785708545 = 119.0
		"01111010", -- (11111110) = -2.0      || 122.40357018327    = 122.0
		"01111101", -- (11111111) = -1.0      || 125.20044652911506 = 125.0

		--	2 => "11111111" , --255
		--	3 => "11010101" ,
		OTHERS => "00000000000"
	);
BEGIN
	---------------
	data_out <= myrom(to_integer(unsigned(address)));
END ARCHITECTURE;