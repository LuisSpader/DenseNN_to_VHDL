LIBRARY ieee;
    USE ieee.std_logic_1164.ALL;
    USE ieee.std_logic_unsigned.ALL;
    USE ieee.numeric_std.ALL;
    USE ieee.math_real.ALL;

    ENTITY  neuron_comb_ReLU_200n_8bit_signed_mul0_v0_add0_v0 IS
        -- GENERIC (
    -- 	input_bit:integer:= 8; output_bit:integer:= 8 ;	 n_input:integer:= 200
        -- );
    PORT (
        clk, rst, update_weights : IN STD_LOGIC;
        x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200: IN signed(7 DOWNTO 0);
    -- 	w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200: IN signed(7 DOWNTO 0);
        bias: IN signed(7 DOWNTO 0) ; -- offset
        ------------------------------------------
        y: OUT signed (7 DOWNTO 0) --output  result
    );
    -- clk, rst,
    -- inputs,
    -- weigths,
    -- bias,
    -- output
    end ENTITY;

    ARCHITECTURE behavior of neuron_comb_ReLU_200n_8bit_signed_mul0_v0_add0_v0 is
    
        COMPONENT MAC_comb_200n_8bit_signed_mul0_v0_add0_v0 IS
        PORT (
            clk, rst : IN STD_LOGIC;
            x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200: IN signed(7 DOWNTO 0);
            w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200: IN signed(7 DOWNTO 0);
            bias: IN signed(7 DOWNTO 0) ; -- offset 
            ------------------------------------------ 
            output: OUT signed(7 DOWNTO 0)
        ); -- clk, rst, inputs, weigths, bias, output
        END COMPONENT;                            
    
    -- # ROM_component
        SIGNAL out_reg_MAC : signed ((7) DOWNTO 0);	--reg da saida do MAC
    
        SIGNAL reg_x1, reg_x2, reg_x3, reg_x4, reg_x5, reg_x6, reg_x7, reg_x8, reg_x9, reg_x10, reg_x11, reg_x12, reg_x13, reg_x14, reg_x15, reg_x16, reg_x17, reg_x18, reg_x19, reg_x20, reg_x21, reg_x22, reg_x23, reg_x24, reg_x25, reg_x26, reg_x27, reg_x28, reg_x29, reg_x30, reg_x31, reg_x32, reg_x33, reg_x34, reg_x35, reg_x36, reg_x37, reg_x38, reg_x39, reg_x40, reg_x41, reg_x42, reg_x43, reg_x44, reg_x45, reg_x46, reg_x47, reg_x48, reg_x49, reg_x50, reg_x51, reg_x52, reg_x53, reg_x54, reg_x55, reg_x56, reg_x57, reg_x58, reg_x59, reg_x60, reg_x61, reg_x62, reg_x63, reg_x64, reg_x65, reg_x66, reg_x67, reg_x68, reg_x69, reg_x70, reg_x71, reg_x72, reg_x73, reg_x74, reg_x75, reg_x76, reg_x77, reg_x78, reg_x79, reg_x80, reg_x81, reg_x82, reg_x83, reg_x84, reg_x85, reg_x86, reg_x87, reg_x88, reg_x89, reg_x90, reg_x91, reg_x92, reg_x93, reg_x94, reg_x95, reg_x96, reg_x97, reg_x98, reg_x99, reg_x100, reg_x101, reg_x102, reg_x103, reg_x104, reg_x105, reg_x106, reg_x107, reg_x108, reg_x109, reg_x110, reg_x111, reg_x112, reg_x113, reg_x114, reg_x115, reg_x116, reg_x117, reg_x118, reg_x119, reg_x120, reg_x121, reg_x122, reg_x123, reg_x124, reg_x125, reg_x126, reg_x127, reg_x128, reg_x129, reg_x130, reg_x131, reg_x132, reg_x133, reg_x134, reg_x135, reg_x136, reg_x137, reg_x138, reg_x139, reg_x140, reg_x141, reg_x142, reg_x143, reg_x144, reg_x145, reg_x146, reg_x147, reg_x148, reg_x149, reg_x150, reg_x151, reg_x152, reg_x153, reg_x154, reg_x155, reg_x156, reg_x157, reg_x158, reg_x159, reg_x160, reg_x161, reg_x162, reg_x163, reg_x164, reg_x165, reg_x166, reg_x167, reg_x168, reg_x169, reg_x170, reg_x171, reg_x172, reg_x173, reg_x174, reg_x175, reg_x176, reg_x177, reg_x178, reg_x179, reg_x180, reg_x181, reg_x182, reg_x183, reg_x184, reg_x185, reg_x186, reg_x187, reg_x188, reg_x189, reg_x190, reg_x191, reg_x192, reg_x193, reg_x194, reg_x195, reg_x196, reg_x197, reg_x198, reg_x199, reg_x200: signed(7 DOWNTO 0); 
        SIGNAL reg_w1, reg_w2, reg_w3, reg_w4, reg_w5, reg_w6, reg_w7, reg_w8, reg_w9, reg_w10, reg_w11, reg_w12, reg_w13, reg_w14, reg_w15, reg_w16, reg_w17, reg_w18, reg_w19, reg_w20, reg_w21, reg_w22, reg_w23, reg_w24, reg_w25, reg_w26, reg_w27, reg_w28, reg_w29, reg_w30, reg_w31, reg_w32, reg_w33, reg_w34, reg_w35, reg_w36, reg_w37, reg_w38, reg_w39, reg_w40, reg_w41, reg_w42, reg_w43, reg_w44, reg_w45, reg_w46, reg_w47, reg_w48, reg_w49, reg_w50, reg_w51, reg_w52, reg_w53, reg_w54, reg_w55, reg_w56, reg_w57, reg_w58, reg_w59, reg_w60, reg_w61, reg_w62, reg_w63, reg_w64, reg_w65, reg_w66, reg_w67, reg_w68, reg_w69, reg_w70, reg_w71, reg_w72, reg_w73, reg_w74, reg_w75, reg_w76, reg_w77, reg_w78, reg_w79, reg_w80, reg_w81, reg_w82, reg_w83, reg_w84, reg_w85, reg_w86, reg_w87, reg_w88, reg_w89, reg_w90, reg_w91, reg_w92, reg_w93, reg_w94, reg_w95, reg_w96, reg_w97, reg_w98, reg_w99, reg_w100, reg_w101, reg_w102, reg_w103, reg_w104, reg_w105, reg_w106, reg_w107, reg_w108, reg_w109, reg_w110, reg_w111, reg_w112, reg_w113, reg_w114, reg_w115, reg_w116, reg_w117, reg_w118, reg_w119, reg_w120, reg_w121, reg_w122, reg_w123, reg_w124, reg_w125, reg_w126, reg_w127, reg_w128, reg_w129, reg_w130, reg_w131, reg_w132, reg_w133, reg_w134, reg_w135, reg_w136, reg_w137, reg_w138, reg_w139, reg_w140, reg_w141, reg_w142, reg_w143, reg_w144, reg_w145, reg_w146, reg_w147, reg_w148, reg_w149, reg_w150, reg_w151, reg_w152, reg_w153, reg_w154, reg_w155, reg_w156, reg_w157, reg_w158, reg_w159, reg_w160, reg_w161, reg_w162, reg_w163, reg_w164, reg_w165, reg_w166, reg_w167, reg_w168, reg_w169, reg_w170, reg_w171, reg_w172, reg_w173, reg_w174, reg_w175, reg_w176, reg_w177, reg_w178, reg_w179, reg_w180, reg_w181, reg_w182, reg_w183, reg_w184, reg_w185, reg_w186, reg_w187, reg_w188, reg_w189, reg_w190, reg_w191, reg_w192, reg_w193, reg_w194, reg_w195, reg_w196, reg_w197, reg_w198, reg_w199, reg_w200: signed(7 DOWNTO 0); 
        SIGNAL reg_bias : signed (7 DOWNTO 0);

    BEGIN
        
        -- MAC ja registra a saida 
	U_MAC : MAC_comb_200n_8bit_signed_mul0_v0_add0_v0 PORT MAP(
            clk, rst, 
	    	reg_x1, reg_x2, reg_x3, reg_x4, reg_x5, reg_x6, reg_x7, reg_x8, reg_x9, reg_x10, reg_x11, reg_x12, reg_x13, reg_x14, reg_x15, reg_x16, reg_x17, reg_x18, reg_x19, reg_x20, reg_x21, reg_x22, reg_x23, reg_x24, reg_x25, reg_x26, reg_x27, reg_x28, reg_x29, reg_x30, reg_x31, reg_x32, reg_x33, reg_x34, reg_x35, reg_x36, reg_x37, reg_x38, reg_x39, reg_x40, reg_x41, reg_x42, reg_x43, reg_x44, reg_x45, reg_x46, reg_x47, reg_x48, reg_x49, reg_x50, reg_x51, reg_x52, reg_x53, reg_x54, reg_x55, reg_x56, reg_x57, reg_x58, reg_x59, reg_x60, reg_x61, reg_x62, reg_x63, reg_x64, reg_x65, reg_x66, reg_x67, reg_x68, reg_x69, reg_x70, reg_x71, reg_x72, reg_x73, reg_x74, reg_x75, reg_x76, reg_x77, reg_x78, reg_x79, reg_x80, reg_x81, reg_x82, reg_x83, reg_x84, reg_x85, reg_x86, reg_x87, reg_x88, reg_x89, reg_x90, reg_x91, reg_x92, reg_x93, reg_x94, reg_x95, reg_x96, reg_x97, reg_x98, reg_x99, reg_x100, reg_x101, reg_x102, reg_x103, reg_x104, reg_x105, reg_x106, reg_x107, reg_x108, reg_x109, reg_x110, reg_x111, reg_x112, reg_x113, reg_x114, reg_x115, reg_x116, reg_x117, reg_x118, reg_x119, reg_x120, reg_x121, reg_x122, reg_x123, reg_x124, reg_x125, reg_x126, reg_x127, reg_x128, reg_x129, reg_x130, reg_x131, reg_x132, reg_x133, reg_x134, reg_x135, reg_x136, reg_x137, reg_x138, reg_x139, reg_x140, reg_x141, reg_x142, reg_x143, reg_x144, reg_x145, reg_x146, reg_x147, reg_x148, reg_x149, reg_x150, reg_x151, reg_x152, reg_x153, reg_x154, reg_x155, reg_x156, reg_x157, reg_x158, reg_x159, reg_x160, reg_x161, reg_x162, reg_x163, reg_x164, reg_x165, reg_x166, reg_x167, reg_x168, reg_x169, reg_x170, reg_x171, reg_x172, reg_x173, reg_x174, reg_x175, reg_x176, reg_x177, reg_x178, reg_x179, reg_x180, reg_x181, reg_x182, reg_x183, reg_x184, reg_x185, reg_x186, reg_x187, reg_x188, reg_x189, reg_x190, reg_x191, reg_x192, reg_x193, reg_x194, reg_x195, reg_x196, reg_x197, reg_x198, reg_x199, reg_x200,
 	   	reg_w1, reg_w2, reg_w3, reg_w4, reg_w5, reg_w6, reg_w7, reg_w8, reg_w9, reg_w10, reg_w11, reg_w12, reg_w13, reg_w14, reg_w15, reg_w16, reg_w17, reg_w18, reg_w19, reg_w20, reg_w21, reg_w22, reg_w23, reg_w24, reg_w25, reg_w26, reg_w27, reg_w28, reg_w29, reg_w30, reg_w31, reg_w32, reg_w33, reg_w34, reg_w35, reg_w36, reg_w37, reg_w38, reg_w39, reg_w40, reg_w41, reg_w42, reg_w43, reg_w44, reg_w45, reg_w46, reg_w47, reg_w48, reg_w49, reg_w50, reg_w51, reg_w52, reg_w53, reg_w54, reg_w55, reg_w56, reg_w57, reg_w58, reg_w59, reg_w60, reg_w61, reg_w62, reg_w63, reg_w64, reg_w65, reg_w66, reg_w67, reg_w68, reg_w69, reg_w70, reg_w71, reg_w72, reg_w73, reg_w74, reg_w75, reg_w76, reg_w77, reg_w78, reg_w79, reg_w80, reg_w81, reg_w82, reg_w83, reg_w84, reg_w85, reg_w86, reg_w87, reg_w88, reg_w89, reg_w90, reg_w91, reg_w92, reg_w93, reg_w94, reg_w95, reg_w96, reg_w97, reg_w98, reg_w99, reg_w100, reg_w101, reg_w102, reg_w103, reg_w104, reg_w105, reg_w106, reg_w107, reg_w108, reg_w109, reg_w110, reg_w111, reg_w112, reg_w113, reg_w114, reg_w115, reg_w116, reg_w117, reg_w118, reg_w119, reg_w120, reg_w121, reg_w122, reg_w123, reg_w124, reg_w125, reg_w126, reg_w127, reg_w128, reg_w129, reg_w130, reg_w131, reg_w132, reg_w133, reg_w134, reg_w135, reg_w136, reg_w137, reg_w138, reg_w139, reg_w140, reg_w141, reg_w142, reg_w143, reg_w144, reg_w145, reg_w146, reg_w147, reg_w148, reg_w149, reg_w150, reg_w151, reg_w152, reg_w153, reg_w154, reg_w155, reg_w156, reg_w157, reg_w158, reg_w159, reg_w160, reg_w161, reg_w162, reg_w163, reg_w164, reg_w165, reg_w166, reg_w167, reg_w168, reg_w169, reg_w170, reg_w171, reg_w172, reg_w173, reg_w174, reg_w175, reg_w176, reg_w177, reg_w178, reg_w179, reg_w180, reg_w181, reg_w182, reg_w183, reg_w184, reg_w185, reg_w186, reg_w187, reg_w188, reg_w189, reg_w190, reg_w191, reg_w192, reg_w193, reg_w194, reg_w195, reg_w196, reg_w197, reg_w198, reg_w199, reg_w200, 
		reg_bias, 
		out_reg_MAC);
        
        PROCESS (clk, rst, update_weights)
        BEGIN
            IF rst = '1' THEN
                                               reg_x1 <= (OTHERS => '0');
                   reg_x2 <= (OTHERS => '0');
                   reg_x3 <= (OTHERS => '0');
                   reg_x4 <= (OTHERS => '0');
                   reg_x5 <= (OTHERS => '0');
                   reg_x6 <= (OTHERS => '0');
                   reg_x7 <= (OTHERS => '0');
                   reg_x8 <= (OTHERS => '0');
                   reg_x9 <= (OTHERS => '0');
                   reg_x10 <= (OTHERS => '0');
                   reg_x11 <= (OTHERS => '0');
                   reg_x12 <= (OTHERS => '0');
                   reg_x13 <= (OTHERS => '0');
                   reg_x14 <= (OTHERS => '0');
                   reg_x15 <= (OTHERS => '0');
                   reg_x16 <= (OTHERS => '0');
                   reg_x17 <= (OTHERS => '0');
                   reg_x18 <= (OTHERS => '0');
                   reg_x19 <= (OTHERS => '0');
                   reg_x20 <= (OTHERS => '0');
                   reg_x21 <= (OTHERS => '0');
                   reg_x22 <= (OTHERS => '0');
                   reg_x23 <= (OTHERS => '0');
                   reg_x24 <= (OTHERS => '0');
                   reg_x25 <= (OTHERS => '0');
                   reg_x26 <= (OTHERS => '0');
                   reg_x27 <= (OTHERS => '0');
                   reg_x28 <= (OTHERS => '0');
                   reg_x29 <= (OTHERS => '0');
                   reg_x30 <= (OTHERS => '0');
                   reg_x31 <= (OTHERS => '0');
                   reg_x32 <= (OTHERS => '0');
                   reg_x33 <= (OTHERS => '0');
                   reg_x34 <= (OTHERS => '0');
                   reg_x35 <= (OTHERS => '0');
                   reg_x36 <= (OTHERS => '0');
                   reg_x37 <= (OTHERS => '0');
                   reg_x38 <= (OTHERS => '0');
                   reg_x39 <= (OTHERS => '0');
                   reg_x40 <= (OTHERS => '0');
                   reg_x41 <= (OTHERS => '0');
                   reg_x42 <= (OTHERS => '0');
                   reg_x43 <= (OTHERS => '0');
                   reg_x44 <= (OTHERS => '0');
                   reg_x45 <= (OTHERS => '0');
                   reg_x46 <= (OTHERS => '0');
                   reg_x47 <= (OTHERS => '0');
                   reg_x48 <= (OTHERS => '0');
                   reg_x49 <= (OTHERS => '0');
                   reg_x50 <= (OTHERS => '0');
                   reg_x51 <= (OTHERS => '0');
                   reg_x52 <= (OTHERS => '0');
                   reg_x53 <= (OTHERS => '0');
                   reg_x54 <= (OTHERS => '0');
                   reg_x55 <= (OTHERS => '0');
                   reg_x56 <= (OTHERS => '0');
                   reg_x57 <= (OTHERS => '0');
                   reg_x58 <= (OTHERS => '0');
                   reg_x59 <= (OTHERS => '0');
                   reg_x60 <= (OTHERS => '0');
                   reg_x61 <= (OTHERS => '0');
                   reg_x62 <= (OTHERS => '0');
                   reg_x63 <= (OTHERS => '0');
                   reg_x64 <= (OTHERS => '0');
                   reg_x65 <= (OTHERS => '0');
                   reg_x66 <= (OTHERS => '0');
                   reg_x67 <= (OTHERS => '0');
                   reg_x68 <= (OTHERS => '0');
                   reg_x69 <= (OTHERS => '0');
                   reg_x70 <= (OTHERS => '0');
                   reg_x71 <= (OTHERS => '0');
                   reg_x72 <= (OTHERS => '0');
                   reg_x73 <= (OTHERS => '0');
                   reg_x74 <= (OTHERS => '0');
                   reg_x75 <= (OTHERS => '0');
                   reg_x76 <= (OTHERS => '0');
                   reg_x77 <= (OTHERS => '0');
                   reg_x78 <= (OTHERS => '0');
                   reg_x79 <= (OTHERS => '0');
                   reg_x80 <= (OTHERS => '0');
                   reg_x81 <= (OTHERS => '0');
                   reg_x82 <= (OTHERS => '0');
                   reg_x83 <= (OTHERS => '0');
                   reg_x84 <= (OTHERS => '0');
                   reg_x85 <= (OTHERS => '0');
                   reg_x86 <= (OTHERS => '0');
                   reg_x87 <= (OTHERS => '0');
                   reg_x88 <= (OTHERS => '0');
                   reg_x89 <= (OTHERS => '0');
                   reg_x90 <= (OTHERS => '0');
                   reg_x91 <= (OTHERS => '0');
                   reg_x92 <= (OTHERS => '0');
                   reg_x93 <= (OTHERS => '0');
                   reg_x94 <= (OTHERS => '0');
                   reg_x95 <= (OTHERS => '0');
                   reg_x96 <= (OTHERS => '0');
                   reg_x97 <= (OTHERS => '0');
                   reg_x98 <= (OTHERS => '0');
                   reg_x99 <= (OTHERS => '0');
                   reg_x100 <= (OTHERS => '0');
                   reg_x101 <= (OTHERS => '0');
                   reg_x102 <= (OTHERS => '0');
                   reg_x103 <= (OTHERS => '0');
                   reg_x104 <= (OTHERS => '0');
                   reg_x105 <= (OTHERS => '0');
                   reg_x106 <= (OTHERS => '0');
                   reg_x107 <= (OTHERS => '0');
                   reg_x108 <= (OTHERS => '0');
                   reg_x109 <= (OTHERS => '0');
                   reg_x110 <= (OTHERS => '0');
                   reg_x111 <= (OTHERS => '0');
                   reg_x112 <= (OTHERS => '0');
                   reg_x113 <= (OTHERS => '0');
                   reg_x114 <= (OTHERS => '0');
                   reg_x115 <= (OTHERS => '0');
                   reg_x116 <= (OTHERS => '0');
                   reg_x117 <= (OTHERS => '0');
                   reg_x118 <= (OTHERS => '0');
                   reg_x119 <= (OTHERS => '0');
                   reg_x120 <= (OTHERS => '0');
                   reg_x121 <= (OTHERS => '0');
                   reg_x122 <= (OTHERS => '0');
                   reg_x123 <= (OTHERS => '0');
                   reg_x124 <= (OTHERS => '0');
                   reg_x125 <= (OTHERS => '0');
                   reg_x126 <= (OTHERS => '0');
                   reg_x127 <= (OTHERS => '0');
                   reg_x128 <= (OTHERS => '0');
                   reg_x129 <= (OTHERS => '0');
                   reg_x130 <= (OTHERS => '0');
                   reg_x131 <= (OTHERS => '0');
                   reg_x132 <= (OTHERS => '0');
                   reg_x133 <= (OTHERS => '0');
                   reg_x134 <= (OTHERS => '0');
                   reg_x135 <= (OTHERS => '0');
                   reg_x136 <= (OTHERS => '0');
                   reg_x137 <= (OTHERS => '0');
                   reg_x138 <= (OTHERS => '0');
                   reg_x139 <= (OTHERS => '0');
                   reg_x140 <= (OTHERS => '0');
                   reg_x141 <= (OTHERS => '0');
                   reg_x142 <= (OTHERS => '0');
                   reg_x143 <= (OTHERS => '0');
                   reg_x144 <= (OTHERS => '0');
                   reg_x145 <= (OTHERS => '0');
                   reg_x146 <= (OTHERS => '0');
                   reg_x147 <= (OTHERS => '0');
                   reg_x148 <= (OTHERS => '0');
                   reg_x149 <= (OTHERS => '0');
                   reg_x150 <= (OTHERS => '0');
                   reg_x151 <= (OTHERS => '0');
                   reg_x152 <= (OTHERS => '0');
                   reg_x153 <= (OTHERS => '0');
                   reg_x154 <= (OTHERS => '0');
                   reg_x155 <= (OTHERS => '0');
                   reg_x156 <= (OTHERS => '0');
                   reg_x157 <= (OTHERS => '0');
                   reg_x158 <= (OTHERS => '0');
                   reg_x159 <= (OTHERS => '0');
                   reg_x160 <= (OTHERS => '0');
                   reg_x161 <= (OTHERS => '0');
                   reg_x162 <= (OTHERS => '0');
                   reg_x163 <= (OTHERS => '0');
                   reg_x164 <= (OTHERS => '0');
                   reg_x165 <= (OTHERS => '0');
                   reg_x166 <= (OTHERS => '0');
                   reg_x167 <= (OTHERS => '0');
                   reg_x168 <= (OTHERS => '0');
                   reg_x169 <= (OTHERS => '0');
                   reg_x170 <= (OTHERS => '0');
                   reg_x171 <= (OTHERS => '0');
                   reg_x172 <= (OTHERS => '0');
                   reg_x173 <= (OTHERS => '0');
                   reg_x174 <= (OTHERS => '0');
                   reg_x175 <= (OTHERS => '0');
                   reg_x176 <= (OTHERS => '0');
                   reg_x177 <= (OTHERS => '0');
                   reg_x178 <= (OTHERS => '0');
                   reg_x179 <= (OTHERS => '0');
                   reg_x180 <= (OTHERS => '0');
                   reg_x181 <= (OTHERS => '0');
                   reg_x182 <= (OTHERS => '0');
                   reg_x183 <= (OTHERS => '0');
                   reg_x184 <= (OTHERS => '0');
                   reg_x185 <= (OTHERS => '0');
                   reg_x186 <= (OTHERS => '0');
                   reg_x187 <= (OTHERS => '0');
                   reg_x188 <= (OTHERS => '0');
                   reg_x189 <= (OTHERS => '0');
                   reg_x190 <= (OTHERS => '0');
                   reg_x191 <= (OTHERS => '0');
                   reg_x192 <= (OTHERS => '0');
                   reg_x193 <= (OTHERS => '0');
                   reg_x194 <= (OTHERS => '0');
                   reg_x195 <= (OTHERS => '0');
                   reg_x196 <= (OTHERS => '0');
                   reg_x197 <= (OTHERS => '0');
                   reg_x198 <= (OTHERS => '0');
                   reg_x199 <= (OTHERS => '0');
                   reg_x200 <= (OTHERS => '0');

                   reg_w1 <= (OTHERS => '0');
                   reg_w2 <= (OTHERS => '0');
                   reg_w3 <= (OTHERS => '0');
                   reg_w4 <= (OTHERS => '0');
                   reg_w5 <= (OTHERS => '0');
                   reg_w6 <= (OTHERS => '0');
                   reg_w7 <= (OTHERS => '0');
                   reg_w8 <= (OTHERS => '0');
                   reg_w9 <= (OTHERS => '0');
                   reg_w10 <= (OTHERS => '0');
                   reg_w11 <= (OTHERS => '0');
                   reg_w12 <= (OTHERS => '0');
                   reg_w13 <= (OTHERS => '0');
                   reg_w14 <= (OTHERS => '0');
                   reg_w15 <= (OTHERS => '0');
                   reg_w16 <= (OTHERS => '0');
                   reg_w17 <= (OTHERS => '0');
                   reg_w18 <= (OTHERS => '0');
                   reg_w19 <= (OTHERS => '0');
                   reg_w20 <= (OTHERS => '0');
                   reg_w21 <= (OTHERS => '0');
                   reg_w22 <= (OTHERS => '0');
                   reg_w23 <= (OTHERS => '0');
                   reg_w24 <= (OTHERS => '0');
                   reg_w25 <= (OTHERS => '0');
                   reg_w26 <= (OTHERS => '0');
                   reg_w27 <= (OTHERS => '0');
                   reg_w28 <= (OTHERS => '0');
                   reg_w29 <= (OTHERS => '0');
                   reg_w30 <= (OTHERS => '0');
                   reg_w31 <= (OTHERS => '0');
                   reg_w32 <= (OTHERS => '0');
                   reg_w33 <= (OTHERS => '0');
                   reg_w34 <= (OTHERS => '0');
                   reg_w35 <= (OTHERS => '0');
                   reg_w36 <= (OTHERS => '0');
                   reg_w37 <= (OTHERS => '0');
                   reg_w38 <= (OTHERS => '0');
                   reg_w39 <= (OTHERS => '0');
                   reg_w40 <= (OTHERS => '0');
                   reg_w41 <= (OTHERS => '0');
                   reg_w42 <= (OTHERS => '0');
                   reg_w43 <= (OTHERS => '0');
                   reg_w44 <= (OTHERS => '0');
                   reg_w45 <= (OTHERS => '0');
                   reg_w46 <= (OTHERS => '0');
                   reg_w47 <= (OTHERS => '0');
                   reg_w48 <= (OTHERS => '0');
                   reg_w49 <= (OTHERS => '0');
                   reg_w50 <= (OTHERS => '0');
                   reg_w51 <= (OTHERS => '0');
                   reg_w52 <= (OTHERS => '0');
                   reg_w53 <= (OTHERS => '0');
                   reg_w54 <= (OTHERS => '0');
                   reg_w55 <= (OTHERS => '0');
                   reg_w56 <= (OTHERS => '0');
                   reg_w57 <= (OTHERS => '0');
                   reg_w58 <= (OTHERS => '0');
                   reg_w59 <= (OTHERS => '0');
                   reg_w60 <= (OTHERS => '0');
                   reg_w61 <= (OTHERS => '0');
                   reg_w62 <= (OTHERS => '0');
                   reg_w63 <= (OTHERS => '0');
                   reg_w64 <= (OTHERS => '0');
                   reg_w65 <= (OTHERS => '0');
                   reg_w66 <= (OTHERS => '0');
                   reg_w67 <= (OTHERS => '0');
                   reg_w68 <= (OTHERS => '0');
                   reg_w69 <= (OTHERS => '0');
                   reg_w70 <= (OTHERS => '0');
                   reg_w71 <= (OTHERS => '0');
                   reg_w72 <= (OTHERS => '0');
                   reg_w73 <= (OTHERS => '0');
                   reg_w74 <= (OTHERS => '0');
                   reg_w75 <= (OTHERS => '0');
                   reg_w76 <= (OTHERS => '0');
                   reg_w77 <= (OTHERS => '0');
                   reg_w78 <= (OTHERS => '0');
                   reg_w79 <= (OTHERS => '0');
                   reg_w80 <= (OTHERS => '0');
                   reg_w81 <= (OTHERS => '0');
                   reg_w82 <= (OTHERS => '0');
                   reg_w83 <= (OTHERS => '0');
                   reg_w84 <= (OTHERS => '0');
                   reg_w85 <= (OTHERS => '0');
                   reg_w86 <= (OTHERS => '0');
                   reg_w87 <= (OTHERS => '0');
                   reg_w88 <= (OTHERS => '0');
                   reg_w89 <= (OTHERS => '0');
                   reg_w90 <= (OTHERS => '0');
                   reg_w91 <= (OTHERS => '0');
                   reg_w92 <= (OTHERS => '0');
                   reg_w93 <= (OTHERS => '0');
                   reg_w94 <= (OTHERS => '0');
                   reg_w95 <= (OTHERS => '0');
                   reg_w96 <= (OTHERS => '0');
                   reg_w97 <= (OTHERS => '0');
                   reg_w98 <= (OTHERS => '0');
                   reg_w99 <= (OTHERS => '0');
                   reg_w100 <= (OTHERS => '0');
                   reg_w101 <= (OTHERS => '0');
                   reg_w102 <= (OTHERS => '0');
                   reg_w103 <= (OTHERS => '0');
                   reg_w104 <= (OTHERS => '0');
                   reg_w105 <= (OTHERS => '0');
                   reg_w106 <= (OTHERS => '0');
                   reg_w107 <= (OTHERS => '0');
                   reg_w108 <= (OTHERS => '0');
                   reg_w109 <= (OTHERS => '0');
                   reg_w110 <= (OTHERS => '0');
                   reg_w111 <= (OTHERS => '0');
                   reg_w112 <= (OTHERS => '0');
                   reg_w113 <= (OTHERS => '0');
                   reg_w114 <= (OTHERS => '0');
                   reg_w115 <= (OTHERS => '0');
                   reg_w116 <= (OTHERS => '0');
                   reg_w117 <= (OTHERS => '0');
                   reg_w118 <= (OTHERS => '0');
                   reg_w119 <= (OTHERS => '0');
                   reg_w120 <= (OTHERS => '0');
                   reg_w121 <= (OTHERS => '0');
                   reg_w122 <= (OTHERS => '0');
                   reg_w123 <= (OTHERS => '0');
                   reg_w124 <= (OTHERS => '0');
                   reg_w125 <= (OTHERS => '0');
                   reg_w126 <= (OTHERS => '0');
                   reg_w127 <= (OTHERS => '0');
                   reg_w128 <= (OTHERS => '0');
                   reg_w129 <= (OTHERS => '0');
                   reg_w130 <= (OTHERS => '0');
                   reg_w131 <= (OTHERS => '0');
                   reg_w132 <= (OTHERS => '0');
                   reg_w133 <= (OTHERS => '0');
                   reg_w134 <= (OTHERS => '0');
                   reg_w135 <= (OTHERS => '0');
                   reg_w136 <= (OTHERS => '0');
                   reg_w137 <= (OTHERS => '0');
                   reg_w138 <= (OTHERS => '0');
                   reg_w139 <= (OTHERS => '0');
                   reg_w140 <= (OTHERS => '0');
                   reg_w141 <= (OTHERS => '0');
                   reg_w142 <= (OTHERS => '0');
                   reg_w143 <= (OTHERS => '0');
                   reg_w144 <= (OTHERS => '0');
                   reg_w145 <= (OTHERS => '0');
                   reg_w146 <= (OTHERS => '0');
                   reg_w147 <= (OTHERS => '0');
                   reg_w148 <= (OTHERS => '0');
                   reg_w149 <= (OTHERS => '0');
                   reg_w150 <= (OTHERS => '0');
                   reg_w151 <= (OTHERS => '0');
                   reg_w152 <= (OTHERS => '0');
                   reg_w153 <= (OTHERS => '0');
                   reg_w154 <= (OTHERS => '0');
                   reg_w155 <= (OTHERS => '0');
                   reg_w156 <= (OTHERS => '0');
                   reg_w157 <= (OTHERS => '0');
                   reg_w158 <= (OTHERS => '0');
                   reg_w159 <= (OTHERS => '0');
                   reg_w160 <= (OTHERS => '0');
                   reg_w161 <= (OTHERS => '0');
                   reg_w162 <= (OTHERS => '0');
                   reg_w163 <= (OTHERS => '0');
                   reg_w164 <= (OTHERS => '0');
                   reg_w165 <= (OTHERS => '0');
                   reg_w166 <= (OTHERS => '0');
                   reg_w167 <= (OTHERS => '0');
                   reg_w168 <= (OTHERS => '0');
                   reg_w169 <= (OTHERS => '0');
                   reg_w170 <= (OTHERS => '0');
                   reg_w171 <= (OTHERS => '0');
                   reg_w172 <= (OTHERS => '0');
                   reg_w173 <= (OTHERS => '0');
                   reg_w174 <= (OTHERS => '0');
                   reg_w175 <= (OTHERS => '0');
                   reg_w176 <= (OTHERS => '0');
                   reg_w177 <= (OTHERS => '0');
                   reg_w178 <= (OTHERS => '0');
                   reg_w179 <= (OTHERS => '0');
                   reg_w180 <= (OTHERS => '0');
                   reg_w181 <= (OTHERS => '0');
                   reg_w182 <= (OTHERS => '0');
                   reg_w183 <= (OTHERS => '0');
                   reg_w184 <= (OTHERS => '0');
                   reg_w185 <= (OTHERS => '0');
                   reg_w186 <= (OTHERS => '0');
                   reg_w187 <= (OTHERS => '0');
                   reg_w188 <= (OTHERS => '0');
                   reg_w189 <= (OTHERS => '0');
                   reg_w190 <= (OTHERS => '0');
                   reg_w191 <= (OTHERS => '0');
                   reg_w192 <= (OTHERS => '0');
                   reg_w193 <= (OTHERS => '0');
                   reg_w194 <= (OTHERS => '0');
                   reg_w195 <= (OTHERS => '0');
                   reg_w196 <= (OTHERS => '0');
                   reg_w197 <= (OTHERS => '0');
                   reg_w198 <= (OTHERS => '0');
                   reg_w199 <= (OTHERS => '0');
                   reg_w200 <= (OTHERS => '0');
                   reg_bias <= (OTHERS => '0');
            ELSIF clk'event AND clk = '1' THEN
        
                IF out_reg_MAC > 0 THEN
                    y <= out_reg_MAC;
                ELSE
                    y <= (OTHERS => '0');
                END IF;
    
                                                   IF update_weights = '0' THEN 
                         reg_x1 <= x1;
                         reg_x2 <= x2;
                         reg_x3 <= x3;
                         reg_x4 <= x4;
                         reg_x5 <= x5;
                         reg_x6 <= x6;
                         reg_x7 <= x7;
                         reg_x8 <= x8;
                         reg_x9 <= x9;
                         reg_x10 <= x10;
                         reg_x11 <= x11;
                         reg_x12 <= x12;
                         reg_x13 <= x13;
                         reg_x14 <= x14;
                         reg_x15 <= x15;
                         reg_x16 <= x16;
                         reg_x17 <= x17;
                         reg_x18 <= x18;
                         reg_x19 <= x19;
                         reg_x20 <= x20;
                         reg_x21 <= x21;
                         reg_x22 <= x22;
                         reg_x23 <= x23;
                         reg_x24 <= x24;
                         reg_x25 <= x25;
                         reg_x26 <= x26;
                         reg_x27 <= x27;
                         reg_x28 <= x28;
                         reg_x29 <= x29;
                         reg_x30 <= x30;
                         reg_x31 <= x31;
                         reg_x32 <= x32;
                         reg_x33 <= x33;
                         reg_x34 <= x34;
                         reg_x35 <= x35;
                         reg_x36 <= x36;
                         reg_x37 <= x37;
                         reg_x38 <= x38;
                         reg_x39 <= x39;
                         reg_x40 <= x40;
                         reg_x41 <= x41;
                         reg_x42 <= x42;
                         reg_x43 <= x43;
                         reg_x44 <= x44;
                         reg_x45 <= x45;
                         reg_x46 <= x46;
                         reg_x47 <= x47;
                         reg_x48 <= x48;
                         reg_x49 <= x49;
                         reg_x50 <= x50;
                         reg_x51 <= x51;
                         reg_x52 <= x52;
                         reg_x53 <= x53;
                         reg_x54 <= x54;
                         reg_x55 <= x55;
                         reg_x56 <= x56;
                         reg_x57 <= x57;
                         reg_x58 <= x58;
                         reg_x59 <= x59;
                         reg_x60 <= x60;
                         reg_x61 <= x61;
                         reg_x62 <= x62;
                         reg_x63 <= x63;
                         reg_x64 <= x64;
                         reg_x65 <= x65;
                         reg_x66 <= x66;
                         reg_x67 <= x67;
                         reg_x68 <= x68;
                         reg_x69 <= x69;
                         reg_x70 <= x70;
                         reg_x71 <= x71;
                         reg_x72 <= x72;
                         reg_x73 <= x73;
                         reg_x74 <= x74;
                         reg_x75 <= x75;
                         reg_x76 <= x76;
                         reg_x77 <= x77;
                         reg_x78 <= x78;
                         reg_x79 <= x79;
                         reg_x80 <= x80;
                         reg_x81 <= x81;
                         reg_x82 <= x82;
                         reg_x83 <= x83;
                         reg_x84 <= x84;
                         reg_x85 <= x85;
                         reg_x86 <= x86;
                         reg_x87 <= x87;
                         reg_x88 <= x88;
                         reg_x89 <= x89;
                         reg_x90 <= x90;
                         reg_x91 <= x91;
                         reg_x92 <= x92;
                         reg_x93 <= x93;
                         reg_x94 <= x94;
                         reg_x95 <= x95;
                         reg_x96 <= x96;
                         reg_x97 <= x97;
                         reg_x98 <= x98;
                         reg_x99 <= x99;
                         reg_x100 <= x100;
                         reg_x101 <= x101;
                         reg_x102 <= x102;
                         reg_x103 <= x103;
                         reg_x104 <= x104;
                         reg_x105 <= x105;
                         reg_x106 <= x106;
                         reg_x107 <= x107;
                         reg_x108 <= x108;
                         reg_x109 <= x109;
                         reg_x110 <= x110;
                         reg_x111 <= x111;
                         reg_x112 <= x112;
                         reg_x113 <= x113;
                         reg_x114 <= x114;
                         reg_x115 <= x115;
                         reg_x116 <= x116;
                         reg_x117 <= x117;
                         reg_x118 <= x118;
                         reg_x119 <= x119;
                         reg_x120 <= x120;
                         reg_x121 <= x121;
                         reg_x122 <= x122;
                         reg_x123 <= x123;
                         reg_x124 <= x124;
                         reg_x125 <= x125;
                         reg_x126 <= x126;
                         reg_x127 <= x127;
                         reg_x128 <= x128;
                         reg_x129 <= x129;
                         reg_x130 <= x130;
                         reg_x131 <= x131;
                         reg_x132 <= x132;
                         reg_x133 <= x133;
                         reg_x134 <= x134;
                         reg_x135 <= x135;
                         reg_x136 <= x136;
                         reg_x137 <= x137;
                         reg_x138 <= x138;
                         reg_x139 <= x139;
                         reg_x140 <= x140;
                         reg_x141 <= x141;
                         reg_x142 <= x142;
                         reg_x143 <= x143;
                         reg_x144 <= x144;
                         reg_x145 <= x145;
                         reg_x146 <= x146;
                         reg_x147 <= x147;
                         reg_x148 <= x148;
                         reg_x149 <= x149;
                         reg_x150 <= x150;
                         reg_x151 <= x151;
                         reg_x152 <= x152;
                         reg_x153 <= x153;
                         reg_x154 <= x154;
                         reg_x155 <= x155;
                         reg_x156 <= x156;
                         reg_x157 <= x157;
                         reg_x158 <= x158;
                         reg_x159 <= x159;
                         reg_x160 <= x160;
                         reg_x161 <= x161;
                         reg_x162 <= x162;
                         reg_x163 <= x163;
                         reg_x164 <= x164;
                         reg_x165 <= x165;
                         reg_x166 <= x166;
                         reg_x167 <= x167;
                         reg_x168 <= x168;
                         reg_x169 <= x169;
                         reg_x170 <= x170;
                         reg_x171 <= x171;
                         reg_x172 <= x172;
                         reg_x173 <= x173;
                         reg_x174 <= x174;
                         reg_x175 <= x175;
                         reg_x176 <= x176;
                         reg_x177 <= x177;
                         reg_x178 <= x178;
                         reg_x179 <= x179;
                         reg_x180 <= x180;
                         reg_x181 <= x181;
                         reg_x182 <= x182;
                         reg_x183 <= x183;
                         reg_x184 <= x184;
                         reg_x185 <= x185;
                         reg_x186 <= x186;
                         reg_x187 <= x187;
                         reg_x188 <= x188;
                         reg_x189 <= x189;
                         reg_x190 <= x190;
                         reg_x191 <= x191;
                         reg_x192 <= x192;
                         reg_x193 <= x193;
                         reg_x194 <= x194;
                         reg_x195 <= x195;
                         reg_x196 <= x196;
                         reg_x197 <= x197;
                         reg_x198 <= x198;
                         reg_x199 <= x199;
                         reg_x200 <= x200;

                       ELSE
                         reg_w1 <= x1;
                         reg_w2 <= x2;
                         reg_w3 <= x3;
                         reg_w4 <= x4;
                         reg_w5 <= x5;
                         reg_w6 <= x6;
                         reg_w7 <= x7;
                         reg_w8 <= x8;
                         reg_w9 <= x9;
                         reg_w10 <= x10;
                         reg_w11 <= x11;
                         reg_w12 <= x12;
                         reg_w13 <= x13;
                         reg_w14 <= x14;
                         reg_w15 <= x15;
                         reg_w16 <= x16;
                         reg_w17 <= x17;
                         reg_w18 <= x18;
                         reg_w19 <= x19;
                         reg_w20 <= x20;
                         reg_w21 <= x21;
                         reg_w22 <= x22;
                         reg_w23 <= x23;
                         reg_w24 <= x24;
                         reg_w25 <= x25;
                         reg_w26 <= x26;
                         reg_w27 <= x27;
                         reg_w28 <= x28;
                         reg_w29 <= x29;
                         reg_w30 <= x30;
                         reg_w31 <= x31;
                         reg_w32 <= x32;
                         reg_w33 <= x33;
                         reg_w34 <= x34;
                         reg_w35 <= x35;
                         reg_w36 <= x36;
                         reg_w37 <= x37;
                         reg_w38 <= x38;
                         reg_w39 <= x39;
                         reg_w40 <= x40;
                         reg_w41 <= x41;
                         reg_w42 <= x42;
                         reg_w43 <= x43;
                         reg_w44 <= x44;
                         reg_w45 <= x45;
                         reg_w46 <= x46;
                         reg_w47 <= x47;
                         reg_w48 <= x48;
                         reg_w49 <= x49;
                         reg_w50 <= x50;
                         reg_w51 <= x51;
                         reg_w52 <= x52;
                         reg_w53 <= x53;
                         reg_w54 <= x54;
                         reg_w55 <= x55;
                         reg_w56 <= x56;
                         reg_w57 <= x57;
                         reg_w58 <= x58;
                         reg_w59 <= x59;
                         reg_w60 <= x60;
                         reg_w61 <= x61;
                         reg_w62 <= x62;
                         reg_w63 <= x63;
                         reg_w64 <= x64;
                         reg_w65 <= x65;
                         reg_w66 <= x66;
                         reg_w67 <= x67;
                         reg_w68 <= x68;
                         reg_w69 <= x69;
                         reg_w70 <= x70;
                         reg_w71 <= x71;
                         reg_w72 <= x72;
                         reg_w73 <= x73;
                         reg_w74 <= x74;
                         reg_w75 <= x75;
                         reg_w76 <= x76;
                         reg_w77 <= x77;
                         reg_w78 <= x78;
                         reg_w79 <= x79;
                         reg_w80 <= x80;
                         reg_w81 <= x81;
                         reg_w82 <= x82;
                         reg_w83 <= x83;
                         reg_w84 <= x84;
                         reg_w85 <= x85;
                         reg_w86 <= x86;
                         reg_w87 <= x87;
                         reg_w88 <= x88;
                         reg_w89 <= x89;
                         reg_w90 <= x90;
                         reg_w91 <= x91;
                         reg_w92 <= x92;
                         reg_w93 <= x93;
                         reg_w94 <= x94;
                         reg_w95 <= x95;
                         reg_w96 <= x96;
                         reg_w97 <= x97;
                         reg_w98 <= x98;
                         reg_w99 <= x99;
                         reg_w100 <= x100;
                         reg_w101 <= x101;
                         reg_w102 <= x102;
                         reg_w103 <= x103;
                         reg_w104 <= x104;
                         reg_w105 <= x105;
                         reg_w106 <= x106;
                         reg_w107 <= x107;
                         reg_w108 <= x108;
                         reg_w109 <= x109;
                         reg_w110 <= x110;
                         reg_w111 <= x111;
                         reg_w112 <= x112;
                         reg_w113 <= x113;
                         reg_w114 <= x114;
                         reg_w115 <= x115;
                         reg_w116 <= x116;
                         reg_w117 <= x117;
                         reg_w118 <= x118;
                         reg_w119 <= x119;
                         reg_w120 <= x120;
                         reg_w121 <= x121;
                         reg_w122 <= x122;
                         reg_w123 <= x123;
                         reg_w124 <= x124;
                         reg_w125 <= x125;
                         reg_w126 <= x126;
                         reg_w127 <= x127;
                         reg_w128 <= x128;
                         reg_w129 <= x129;
                         reg_w130 <= x130;
                         reg_w131 <= x131;
                         reg_w132 <= x132;
                         reg_w133 <= x133;
                         reg_w134 <= x134;
                         reg_w135 <= x135;
                         reg_w136 <= x136;
                         reg_w137 <= x137;
                         reg_w138 <= x138;
                         reg_w139 <= x139;
                         reg_w140 <= x140;
                         reg_w141 <= x141;
                         reg_w142 <= x142;
                         reg_w143 <= x143;
                         reg_w144 <= x144;
                         reg_w145 <= x145;
                         reg_w146 <= x146;
                         reg_w147 <= x147;
                         reg_w148 <= x148;
                         reg_w149 <= x149;
                         reg_w150 <= x150;
                         reg_w151 <= x151;
                         reg_w152 <= x152;
                         reg_w153 <= x153;
                         reg_w154 <= x154;
                         reg_w155 <= x155;
                         reg_w156 <= x156;
                         reg_w157 <= x157;
                         reg_w158 <= x158;
                         reg_w159 <= x159;
                         reg_w160 <= x160;
                         reg_w161 <= x161;
                         reg_w162 <= x162;
                         reg_w163 <= x163;
                         reg_w164 <= x164;
                         reg_w165 <= x165;
                         reg_w166 <= x166;
                         reg_w167 <= x167;
                         reg_w168 <= x168;
                         reg_w169 <= x169;
                         reg_w170 <= x170;
                         reg_w171 <= x171;
                         reg_w172 <= x172;
                         reg_w173 <= x173;
                         reg_w174 <= x174;
                         reg_w175 <= x175;
                         reg_w176 <= x176;
                         reg_w177 <= x177;
                         reg_w178 <= x178;
                         reg_w179 <= x179;
                         reg_w180 <= x180;
                         reg_w181 <= x181;
                         reg_w182 <= x182;
                         reg_w183 <= x183;
                         reg_w184 <= x184;
                         reg_w185 <= x185;
                         reg_w186 <= x186;
                         reg_w187 <= x187;
                         reg_w188 <= x188;
                         reg_w189 <= x189;
                         reg_w190 <= x190;
                         reg_w191 <= x191;
                         reg_w192 <= x192;
                         reg_w193 <= x193;
                         reg_w194 <= x194;
                         reg_w195 <= x195;
                         reg_w196 <= x196;
                         reg_w197 <= x197;
                         reg_w198 <= x198;
                         reg_w199 <= x199;
                         reg_w200 <= x200;

                       END IF;
                       reg_bias <= bias;
            END IF;
        END PROCESS;
    
    END behavior;