LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada0_ReLU_10neuron_8bits_200n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c0_n0_bias, c0_n1_bias, c0_n2_bias, c0_n3_bias, c0_n4_bias, c0_n5_bias, c0_n6_bias, c0_n7_bias, c0_n8_bias, c0_n9_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, c0_n0_w1, c0_n0_w2, c0_n0_w3, c0_n0_w4, c0_n0_w5, c0_n0_w6, c0_n0_w7, c0_n0_w8, c0_n0_w9, c0_n0_w10, c0_n0_w11, c0_n0_w12, c0_n0_w13, c0_n0_w14, c0_n0_w15, c0_n0_w16, c0_n0_w17, c0_n0_w18, c0_n0_w19, c0_n0_w20, c0_n0_w21, c0_n0_w22, c0_n0_w23, c0_n0_w24, c0_n0_w25, c0_n0_w26, c0_n0_w27, c0_n0_w28, c0_n0_w29, c0_n0_w30, c0_n0_w31, c0_n0_w32, c0_n0_w33, c0_n0_w34, c0_n0_w35, c0_n0_w36, c0_n0_w37, c0_n0_w38, c0_n0_w39, c0_n0_w40, c0_n0_w41, c0_n0_w42, c0_n0_w43, c0_n0_w44, c0_n0_w45, c0_n0_w46, c0_n0_w47, c0_n0_w48, c0_n0_w49, c0_n0_w50, c0_n0_w51, c0_n0_w52, c0_n0_w53, c0_n0_w54, c0_n0_w55, c0_n0_w56, c0_n0_w57, c0_n0_w58, c0_n0_w59, c0_n0_w60, c0_n0_w61, c0_n0_w62, c0_n0_w63, c0_n0_w64, c0_n0_w65, c0_n0_w66, c0_n0_w67, c0_n0_w68, c0_n0_w69, c0_n0_w70, c0_n0_w71, c0_n0_w72, c0_n0_w73, c0_n0_w74, c0_n0_w75, c0_n0_w76, c0_n0_w77, c0_n0_w78, c0_n0_w79, c0_n0_w80, c0_n0_w81, c0_n0_w82, c0_n0_w83, c0_n0_w84, c0_n0_w85, c0_n0_w86, c0_n0_w87, c0_n0_w88, c0_n0_w89, c0_n0_w90, c0_n0_w91, c0_n0_w92, c0_n0_w93, c0_n0_w94, c0_n0_w95, c0_n0_w96, c0_n0_w97, c0_n0_w98, c0_n0_w99, c0_n0_w100, c0_n0_w101, c0_n0_w102, c0_n0_w103, c0_n0_w104, c0_n0_w105, c0_n0_w106, c0_n0_w107, c0_n0_w108, c0_n0_w109, c0_n0_w110, c0_n0_w111, c0_n0_w112, c0_n0_w113, c0_n0_w114, c0_n0_w115, c0_n0_w116, c0_n0_w117, c0_n0_w118, c0_n0_w119, c0_n0_w120, c0_n0_w121, c0_n0_w122, c0_n0_w123, c0_n0_w124, c0_n0_w125, c0_n0_w126, c0_n0_w127, c0_n0_w128, c0_n0_w129, c0_n0_w130, c0_n0_w131, c0_n0_w132, c0_n0_w133, c0_n0_w134, c0_n0_w135, c0_n0_w136, c0_n0_w137, c0_n0_w138, c0_n0_w139, c0_n0_w140, c0_n0_w141, c0_n0_w142, c0_n0_w143, c0_n0_w144, c0_n0_w145, c0_n0_w146, c0_n0_w147, c0_n0_w148, c0_n0_w149, c0_n0_w150, c0_n0_w151, c0_n0_w152, c0_n0_w153, c0_n0_w154, c0_n0_w155, c0_n0_w156, c0_n0_w157, c0_n0_w158, c0_n0_w159, c0_n0_w160, c0_n0_w161, c0_n0_w162, c0_n0_w163, c0_n0_w164, c0_n0_w165, c0_n0_w166, c0_n0_w167, c0_n0_w168, c0_n0_w169, c0_n0_w170, c0_n0_w171, c0_n0_w172, c0_n0_w173, c0_n0_w174, c0_n0_w175, c0_n0_w176, c0_n0_w177, c0_n0_w178, c0_n0_w179, c0_n0_w180, c0_n0_w181, c0_n0_w182, c0_n0_w183, c0_n0_w184, c0_n0_w185, c0_n0_w186, c0_n0_w187, c0_n0_w188, c0_n0_w189, c0_n0_w190, c0_n0_w191, c0_n0_w192, c0_n0_w193, c0_n0_w194, c0_n0_w195, c0_n0_w196, c0_n0_w197, c0_n0_w198, c0_n0_w199, c0_n0_w200, c0_n1_w1, c0_n1_w2, c0_n1_w3, c0_n1_w4, c0_n1_w5, c0_n1_w6, c0_n1_w7, c0_n1_w8, c0_n1_w9, c0_n1_w10, c0_n1_w11, c0_n1_w12, c0_n1_w13, c0_n1_w14, c0_n1_w15, c0_n1_w16, c0_n1_w17, c0_n1_w18, c0_n1_w19, c0_n1_w20, c0_n1_w21, c0_n1_w22, c0_n1_w23, c0_n1_w24, c0_n1_w25, c0_n1_w26, c0_n1_w27, c0_n1_w28, c0_n1_w29, c0_n1_w30, c0_n1_w31, c0_n1_w32, c0_n1_w33, c0_n1_w34, c0_n1_w35, c0_n1_w36, c0_n1_w37, c0_n1_w38, c0_n1_w39, c0_n1_w40, c0_n1_w41, c0_n1_w42, c0_n1_w43, c0_n1_w44, c0_n1_w45, c0_n1_w46, c0_n1_w47, c0_n1_w48, c0_n1_w49, c0_n1_w50, c0_n1_w51, c0_n1_w52, c0_n1_w53, c0_n1_w54, c0_n1_w55, c0_n1_w56, c0_n1_w57, c0_n1_w58, c0_n1_w59, c0_n1_w60, c0_n1_w61, c0_n1_w62, c0_n1_w63, c0_n1_w64, c0_n1_w65, c0_n1_w66, c0_n1_w67, c0_n1_w68, c0_n1_w69, c0_n1_w70, c0_n1_w71, c0_n1_w72, c0_n1_w73, c0_n1_w74, c0_n1_w75, c0_n1_w76, c0_n1_w77, c0_n1_w78, c0_n1_w79, c0_n1_w80, c0_n1_w81, c0_n1_w82, c0_n1_w83, c0_n1_w84, c0_n1_w85, c0_n1_w86, c0_n1_w87, c0_n1_w88, c0_n1_w89, c0_n1_w90, c0_n1_w91, c0_n1_w92, c0_n1_w93, c0_n1_w94, c0_n1_w95, c0_n1_w96, c0_n1_w97, c0_n1_w98, c0_n1_w99, c0_n1_w100, c0_n1_w101, c0_n1_w102, c0_n1_w103, c0_n1_w104, c0_n1_w105, c0_n1_w106, c0_n1_w107, c0_n1_w108, c0_n1_w109, c0_n1_w110, c0_n1_w111, c0_n1_w112, c0_n1_w113, c0_n1_w114, c0_n1_w115, c0_n1_w116, c0_n1_w117, c0_n1_w118, c0_n1_w119, c0_n1_w120, c0_n1_w121, c0_n1_w122, c0_n1_w123, c0_n1_w124, c0_n1_w125, c0_n1_w126, c0_n1_w127, c0_n1_w128, c0_n1_w129, c0_n1_w130, c0_n1_w131, c0_n1_w132, c0_n1_w133, c0_n1_w134, c0_n1_w135, c0_n1_w136, c0_n1_w137, c0_n1_w138, c0_n1_w139, c0_n1_w140, c0_n1_w141, c0_n1_w142, c0_n1_w143, c0_n1_w144, c0_n1_w145, c0_n1_w146, c0_n1_w147, c0_n1_w148, c0_n1_w149, c0_n1_w150, c0_n1_w151, c0_n1_w152, c0_n1_w153, c0_n1_w154, c0_n1_w155, c0_n1_w156, c0_n1_w157, c0_n1_w158, c0_n1_w159, c0_n1_w160, c0_n1_w161, c0_n1_w162, c0_n1_w163, c0_n1_w164, c0_n1_w165, c0_n1_w166, c0_n1_w167, c0_n1_w168, c0_n1_w169, c0_n1_w170, c0_n1_w171, c0_n1_w172, c0_n1_w173, c0_n1_w174, c0_n1_w175, c0_n1_w176, c0_n1_w177, c0_n1_w178, c0_n1_w179, c0_n1_w180, c0_n1_w181, c0_n1_w182, c0_n1_w183, c0_n1_w184, c0_n1_w185, c0_n1_w186, c0_n1_w187, c0_n1_w188, c0_n1_w189, c0_n1_w190, c0_n1_w191, c0_n1_w192, c0_n1_w193, c0_n1_w194, c0_n1_w195, c0_n1_w196, c0_n1_w197, c0_n1_w198, c0_n1_w199, c0_n1_w200, c0_n2_w1, c0_n2_w2, c0_n2_w3, c0_n2_w4, c0_n2_w5, c0_n2_w6, c0_n2_w7, c0_n2_w8, c0_n2_w9, c0_n2_w10, c0_n2_w11, c0_n2_w12, c0_n2_w13, c0_n2_w14, c0_n2_w15, c0_n2_w16, c0_n2_w17, c0_n2_w18, c0_n2_w19, c0_n2_w20, c0_n2_w21, c0_n2_w22, c0_n2_w23, c0_n2_w24, c0_n2_w25, c0_n2_w26, c0_n2_w27, c0_n2_w28, c0_n2_w29, c0_n2_w30, c0_n2_w31, c0_n2_w32, c0_n2_w33, c0_n2_w34, c0_n2_w35, c0_n2_w36, c0_n2_w37, c0_n2_w38, c0_n2_w39, c0_n2_w40, c0_n2_w41, c0_n2_w42, c0_n2_w43, c0_n2_w44, c0_n2_w45, c0_n2_w46, c0_n2_w47, c0_n2_w48, c0_n2_w49, c0_n2_w50, c0_n2_w51, c0_n2_w52, c0_n2_w53, c0_n2_w54, c0_n2_w55, c0_n2_w56, c0_n2_w57, c0_n2_w58, c0_n2_w59, c0_n2_w60, c0_n2_w61, c0_n2_w62, c0_n2_w63, c0_n2_w64, c0_n2_w65, c0_n2_w66, c0_n2_w67, c0_n2_w68, c0_n2_w69, c0_n2_w70, c0_n2_w71, c0_n2_w72, c0_n2_w73, c0_n2_w74, c0_n2_w75, c0_n2_w76, c0_n2_w77, c0_n2_w78, c0_n2_w79, c0_n2_w80, c0_n2_w81, c0_n2_w82, c0_n2_w83, c0_n2_w84, c0_n2_w85, c0_n2_w86, c0_n2_w87, c0_n2_w88, c0_n2_w89, c0_n2_w90, c0_n2_w91, c0_n2_w92, c0_n2_w93, c0_n2_w94, c0_n2_w95, c0_n2_w96, c0_n2_w97, c0_n2_w98, c0_n2_w99, c0_n2_w100, c0_n2_w101, c0_n2_w102, c0_n2_w103, c0_n2_w104, c0_n2_w105, c0_n2_w106, c0_n2_w107, c0_n2_w108, c0_n2_w109, c0_n2_w110, c0_n2_w111, c0_n2_w112, c0_n2_w113, c0_n2_w114, c0_n2_w115, c0_n2_w116, c0_n2_w117, c0_n2_w118, c0_n2_w119, c0_n2_w120, c0_n2_w121, c0_n2_w122, c0_n2_w123, c0_n2_w124, c0_n2_w125, c0_n2_w126, c0_n2_w127, c0_n2_w128, c0_n2_w129, c0_n2_w130, c0_n2_w131, c0_n2_w132, c0_n2_w133, c0_n2_w134, c0_n2_w135, c0_n2_w136, c0_n2_w137, c0_n2_w138, c0_n2_w139, c0_n2_w140, c0_n2_w141, c0_n2_w142, c0_n2_w143, c0_n2_w144, c0_n2_w145, c0_n2_w146, c0_n2_w147, c0_n2_w148, c0_n2_w149, c0_n2_w150, c0_n2_w151, c0_n2_w152, c0_n2_w153, c0_n2_w154, c0_n2_w155, c0_n2_w156, c0_n2_w157, c0_n2_w158, c0_n2_w159, c0_n2_w160, c0_n2_w161, c0_n2_w162, c0_n2_w163, c0_n2_w164, c0_n2_w165, c0_n2_w166, c0_n2_w167, c0_n2_w168, c0_n2_w169, c0_n2_w170, c0_n2_w171, c0_n2_w172, c0_n2_w173, c0_n2_w174, c0_n2_w175, c0_n2_w176, c0_n2_w177, c0_n2_w178, c0_n2_w179, c0_n2_w180, c0_n2_w181, c0_n2_w182, c0_n2_w183, c0_n2_w184, c0_n2_w185, c0_n2_w186, c0_n2_w187, c0_n2_w188, c0_n2_w189, c0_n2_w190, c0_n2_w191, c0_n2_w192, c0_n2_w193, c0_n2_w194, c0_n2_w195, c0_n2_w196, c0_n2_w197, c0_n2_w198, c0_n2_w199, c0_n2_w200, c0_n3_w1, c0_n3_w2, c0_n3_w3, c0_n3_w4, c0_n3_w5, c0_n3_w6, c0_n3_w7, c0_n3_w8, c0_n3_w9, c0_n3_w10, c0_n3_w11, c0_n3_w12, c0_n3_w13, c0_n3_w14, c0_n3_w15, c0_n3_w16, c0_n3_w17, c0_n3_w18, c0_n3_w19, c0_n3_w20, c0_n3_w21, c0_n3_w22, c0_n3_w23, c0_n3_w24, c0_n3_w25, c0_n3_w26, c0_n3_w27, c0_n3_w28, c0_n3_w29, c0_n3_w30, c0_n3_w31, c0_n3_w32, c0_n3_w33, c0_n3_w34, c0_n3_w35, c0_n3_w36, c0_n3_w37, c0_n3_w38, c0_n3_w39, c0_n3_w40, c0_n3_w41, c0_n3_w42, c0_n3_w43, c0_n3_w44, c0_n3_w45, c0_n3_w46, c0_n3_w47, c0_n3_w48, c0_n3_w49, c0_n3_w50, c0_n3_w51, c0_n3_w52, c0_n3_w53, c0_n3_w54, c0_n3_w55, c0_n3_w56, c0_n3_w57, c0_n3_w58, c0_n3_w59, c0_n3_w60, c0_n3_w61, c0_n3_w62, c0_n3_w63, c0_n3_w64, c0_n3_w65, c0_n3_w66, c0_n3_w67, c0_n3_w68, c0_n3_w69, c0_n3_w70, c0_n3_w71, c0_n3_w72, c0_n3_w73, c0_n3_w74, c0_n3_w75, c0_n3_w76, c0_n3_w77, c0_n3_w78, c0_n3_w79, c0_n3_w80, c0_n3_w81, c0_n3_w82, c0_n3_w83, c0_n3_w84, c0_n3_w85, c0_n3_w86, c0_n3_w87, c0_n3_w88, c0_n3_w89, c0_n3_w90, c0_n3_w91, c0_n3_w92, c0_n3_w93, c0_n3_w94, c0_n3_w95, c0_n3_w96, c0_n3_w97, c0_n3_w98, c0_n3_w99, c0_n3_w100, c0_n3_w101, c0_n3_w102, c0_n3_w103, c0_n3_w104, c0_n3_w105, c0_n3_w106, c0_n3_w107, c0_n3_w108, c0_n3_w109, c0_n3_w110, c0_n3_w111, c0_n3_w112, c0_n3_w113, c0_n3_w114, c0_n3_w115, c0_n3_w116, c0_n3_w117, c0_n3_w118, c0_n3_w119, c0_n3_w120, c0_n3_w121, c0_n3_w122, c0_n3_w123, c0_n3_w124, c0_n3_w125, c0_n3_w126, c0_n3_w127, c0_n3_w128, c0_n3_w129, c0_n3_w130, c0_n3_w131, c0_n3_w132, c0_n3_w133, c0_n3_w134, c0_n3_w135, c0_n3_w136, c0_n3_w137, c0_n3_w138, c0_n3_w139, c0_n3_w140, c0_n3_w141, c0_n3_w142, c0_n3_w143, c0_n3_w144, c0_n3_w145, c0_n3_w146, c0_n3_w147, c0_n3_w148, c0_n3_w149, c0_n3_w150, c0_n3_w151, c0_n3_w152, c0_n3_w153, c0_n3_w154, c0_n3_w155, c0_n3_w156, c0_n3_w157, c0_n3_w158, c0_n3_w159, c0_n3_w160, c0_n3_w161, c0_n3_w162, c0_n3_w163, c0_n3_w164, c0_n3_w165, c0_n3_w166, c0_n3_w167, c0_n3_w168, c0_n3_w169, c0_n3_w170, c0_n3_w171, c0_n3_w172, c0_n3_w173, c0_n3_w174, c0_n3_w175, c0_n3_w176, c0_n3_w177, c0_n3_w178, c0_n3_w179, c0_n3_w180, c0_n3_w181, c0_n3_w182, c0_n3_w183, c0_n3_w184, c0_n3_w185, c0_n3_w186, c0_n3_w187, c0_n3_w188, c0_n3_w189, c0_n3_w190, c0_n3_w191, c0_n3_w192, c0_n3_w193, c0_n3_w194, c0_n3_w195, c0_n3_w196, c0_n3_w197, c0_n3_w198, c0_n3_w199, c0_n3_w200, c0_n4_w1, c0_n4_w2, c0_n4_w3, c0_n4_w4, c0_n4_w5, c0_n4_w6, c0_n4_w7, c0_n4_w8, c0_n4_w9, c0_n4_w10, c0_n4_w11, c0_n4_w12, c0_n4_w13, c0_n4_w14, c0_n4_w15, c0_n4_w16, c0_n4_w17, c0_n4_w18, c0_n4_w19, c0_n4_w20, c0_n4_w21, c0_n4_w22, c0_n4_w23, c0_n4_w24, c0_n4_w25, c0_n4_w26, c0_n4_w27, c0_n4_w28, c0_n4_w29, c0_n4_w30, c0_n4_w31, c0_n4_w32, c0_n4_w33, c0_n4_w34, c0_n4_w35, c0_n4_w36, c0_n4_w37, c0_n4_w38, c0_n4_w39, c0_n4_w40, c0_n4_w41, c0_n4_w42, c0_n4_w43, c0_n4_w44, c0_n4_w45, c0_n4_w46, c0_n4_w47, c0_n4_w48, c0_n4_w49, c0_n4_w50, c0_n4_w51, c0_n4_w52, c0_n4_w53, c0_n4_w54, c0_n4_w55, c0_n4_w56, c0_n4_w57, c0_n4_w58, c0_n4_w59, c0_n4_w60, c0_n4_w61, c0_n4_w62, c0_n4_w63, c0_n4_w64, c0_n4_w65, c0_n4_w66, c0_n4_w67, c0_n4_w68, c0_n4_w69, c0_n4_w70, c0_n4_w71, c0_n4_w72, c0_n4_w73, c0_n4_w74, c0_n4_w75, c0_n4_w76, c0_n4_w77, c0_n4_w78, c0_n4_w79, c0_n4_w80, c0_n4_w81, c0_n4_w82, c0_n4_w83, c0_n4_w84, c0_n4_w85, c0_n4_w86, c0_n4_w87, c0_n4_w88, c0_n4_w89, c0_n4_w90, c0_n4_w91, c0_n4_w92, c0_n4_w93, c0_n4_w94, c0_n4_w95, c0_n4_w96, c0_n4_w97, c0_n4_w98, c0_n4_w99, c0_n4_w100, c0_n4_w101, c0_n4_w102, c0_n4_w103, c0_n4_w104, c0_n4_w105, c0_n4_w106, c0_n4_w107, c0_n4_w108, c0_n4_w109, c0_n4_w110, c0_n4_w111, c0_n4_w112, c0_n4_w113, c0_n4_w114, c0_n4_w115, c0_n4_w116, c0_n4_w117, c0_n4_w118, c0_n4_w119, c0_n4_w120, c0_n4_w121, c0_n4_w122, c0_n4_w123, c0_n4_w124, c0_n4_w125, c0_n4_w126, c0_n4_w127, c0_n4_w128, c0_n4_w129, c0_n4_w130, c0_n4_w131, c0_n4_w132, c0_n4_w133, c0_n4_w134, c0_n4_w135, c0_n4_w136, c0_n4_w137, c0_n4_w138, c0_n4_w139, c0_n4_w140, c0_n4_w141, c0_n4_w142, c0_n4_w143, c0_n4_w144, c0_n4_w145, c0_n4_w146, c0_n4_w147, c0_n4_w148, c0_n4_w149, c0_n4_w150, c0_n4_w151, c0_n4_w152, c0_n4_w153, c0_n4_w154, c0_n4_w155, c0_n4_w156, c0_n4_w157, c0_n4_w158, c0_n4_w159, c0_n4_w160, c0_n4_w161, c0_n4_w162, c0_n4_w163, c0_n4_w164, c0_n4_w165, c0_n4_w166, c0_n4_w167, c0_n4_w168, c0_n4_w169, c0_n4_w170, c0_n4_w171, c0_n4_w172, c0_n4_w173, c0_n4_w174, c0_n4_w175, c0_n4_w176, c0_n4_w177, c0_n4_w178, c0_n4_w179, c0_n4_w180, c0_n4_w181, c0_n4_w182, c0_n4_w183, c0_n4_w184, c0_n4_w185, c0_n4_w186, c0_n4_w187, c0_n4_w188, c0_n4_w189, c0_n4_w190, c0_n4_w191, c0_n4_w192, c0_n4_w193, c0_n4_w194, c0_n4_w195, c0_n4_w196, c0_n4_w197, c0_n4_w198, c0_n4_w199, c0_n4_w200, c0_n5_w1, c0_n5_w2, c0_n5_w3, c0_n5_w4, c0_n5_w5, c0_n5_w6, c0_n5_w7, c0_n5_w8, c0_n5_w9, c0_n5_w10, c0_n5_w11, c0_n5_w12, c0_n5_w13, c0_n5_w14, c0_n5_w15, c0_n5_w16, c0_n5_w17, c0_n5_w18, c0_n5_w19, c0_n5_w20, c0_n5_w21, c0_n5_w22, c0_n5_w23, c0_n5_w24, c0_n5_w25, c0_n5_w26, c0_n5_w27, c0_n5_w28, c0_n5_w29, c0_n5_w30, c0_n5_w31, c0_n5_w32, c0_n5_w33, c0_n5_w34, c0_n5_w35, c0_n5_w36, c0_n5_w37, c0_n5_w38, c0_n5_w39, c0_n5_w40, c0_n5_w41, c0_n5_w42, c0_n5_w43, c0_n5_w44, c0_n5_w45, c0_n5_w46, c0_n5_w47, c0_n5_w48, c0_n5_w49, c0_n5_w50, c0_n5_w51, c0_n5_w52, c0_n5_w53, c0_n5_w54, c0_n5_w55, c0_n5_w56, c0_n5_w57, c0_n5_w58, c0_n5_w59, c0_n5_w60, c0_n5_w61, c0_n5_w62, c0_n5_w63, c0_n5_w64, c0_n5_w65, c0_n5_w66, c0_n5_w67, c0_n5_w68, c0_n5_w69, c0_n5_w70, c0_n5_w71, c0_n5_w72, c0_n5_w73, c0_n5_w74, c0_n5_w75, c0_n5_w76, c0_n5_w77, c0_n5_w78, c0_n5_w79, c0_n5_w80, c0_n5_w81, c0_n5_w82, c0_n5_w83, c0_n5_w84, c0_n5_w85, c0_n5_w86, c0_n5_w87, c0_n5_w88, c0_n5_w89, c0_n5_w90, c0_n5_w91, c0_n5_w92, c0_n5_w93, c0_n5_w94, c0_n5_w95, c0_n5_w96, c0_n5_w97, c0_n5_w98, c0_n5_w99, c0_n5_w100, c0_n5_w101, c0_n5_w102, c0_n5_w103, c0_n5_w104, c0_n5_w105, c0_n5_w106, c0_n5_w107, c0_n5_w108, c0_n5_w109, c0_n5_w110, c0_n5_w111, c0_n5_w112, c0_n5_w113, c0_n5_w114, c0_n5_w115, c0_n5_w116, c0_n5_w117, c0_n5_w118, c0_n5_w119, c0_n5_w120, c0_n5_w121, c0_n5_w122, c0_n5_w123, c0_n5_w124, c0_n5_w125, c0_n5_w126, c0_n5_w127, c0_n5_w128, c0_n5_w129, c0_n5_w130, c0_n5_w131, c0_n5_w132, c0_n5_w133, c0_n5_w134, c0_n5_w135, c0_n5_w136, c0_n5_w137, c0_n5_w138, c0_n5_w139, c0_n5_w140, c0_n5_w141, c0_n5_w142, c0_n5_w143, c0_n5_w144, c0_n5_w145, c0_n5_w146, c0_n5_w147, c0_n5_w148, c0_n5_w149, c0_n5_w150, c0_n5_w151, c0_n5_w152, c0_n5_w153, c0_n5_w154, c0_n5_w155, c0_n5_w156, c0_n5_w157, c0_n5_w158, c0_n5_w159, c0_n5_w160, c0_n5_w161, c0_n5_w162, c0_n5_w163, c0_n5_w164, c0_n5_w165, c0_n5_w166, c0_n5_w167, c0_n5_w168, c0_n5_w169, c0_n5_w170, c0_n5_w171, c0_n5_w172, c0_n5_w173, c0_n5_w174, c0_n5_w175, c0_n5_w176, c0_n5_w177, c0_n5_w178, c0_n5_w179, c0_n5_w180, c0_n5_w181, c0_n5_w182, c0_n5_w183, c0_n5_w184, c0_n5_w185, c0_n5_w186, c0_n5_w187, c0_n5_w188, c0_n5_w189, c0_n5_w190, c0_n5_w191, c0_n5_w192, c0_n5_w193, c0_n5_w194, c0_n5_w195, c0_n5_w196, c0_n5_w197, c0_n5_w198, c0_n5_w199, c0_n5_w200, c0_n6_w1, c0_n6_w2, c0_n6_w3, c0_n6_w4, c0_n6_w5, c0_n6_w6, c0_n6_w7, c0_n6_w8, c0_n6_w9, c0_n6_w10, c0_n6_w11, c0_n6_w12, c0_n6_w13, c0_n6_w14, c0_n6_w15, c0_n6_w16, c0_n6_w17, c0_n6_w18, c0_n6_w19, c0_n6_w20, c0_n6_w21, c0_n6_w22, c0_n6_w23, c0_n6_w24, c0_n6_w25, c0_n6_w26, c0_n6_w27, c0_n6_w28, c0_n6_w29, c0_n6_w30, c0_n6_w31, c0_n6_w32, c0_n6_w33, c0_n6_w34, c0_n6_w35, c0_n6_w36, c0_n6_w37, c0_n6_w38, c0_n6_w39, c0_n6_w40, c0_n6_w41, c0_n6_w42, c0_n6_w43, c0_n6_w44, c0_n6_w45, c0_n6_w46, c0_n6_w47, c0_n6_w48, c0_n6_w49, c0_n6_w50, c0_n6_w51, c0_n6_w52, c0_n6_w53, c0_n6_w54, c0_n6_w55, c0_n6_w56, c0_n6_w57, c0_n6_w58, c0_n6_w59, c0_n6_w60, c0_n6_w61, c0_n6_w62, c0_n6_w63, c0_n6_w64, c0_n6_w65, c0_n6_w66, c0_n6_w67, c0_n6_w68, c0_n6_w69, c0_n6_w70, c0_n6_w71, c0_n6_w72, c0_n6_w73, c0_n6_w74, c0_n6_w75, c0_n6_w76, c0_n6_w77, c0_n6_w78, c0_n6_w79, c0_n6_w80, c0_n6_w81, c0_n6_w82, c0_n6_w83, c0_n6_w84, c0_n6_w85, c0_n6_w86, c0_n6_w87, c0_n6_w88, c0_n6_w89, c0_n6_w90, c0_n6_w91, c0_n6_w92, c0_n6_w93, c0_n6_w94, c0_n6_w95, c0_n6_w96, c0_n6_w97, c0_n6_w98, c0_n6_w99, c0_n6_w100, c0_n6_w101, c0_n6_w102, c0_n6_w103, c0_n6_w104, c0_n6_w105, c0_n6_w106, c0_n6_w107, c0_n6_w108, c0_n6_w109, c0_n6_w110, c0_n6_w111, c0_n6_w112, c0_n6_w113, c0_n6_w114, c0_n6_w115, c0_n6_w116, c0_n6_w117, c0_n6_w118, c0_n6_w119, c0_n6_w120, c0_n6_w121, c0_n6_w122, c0_n6_w123, c0_n6_w124, c0_n6_w125, c0_n6_w126, c0_n6_w127, c0_n6_w128, c0_n6_w129, c0_n6_w130, c0_n6_w131, c0_n6_w132, c0_n6_w133, c0_n6_w134, c0_n6_w135, c0_n6_w136, c0_n6_w137, c0_n6_w138, c0_n6_w139, c0_n6_w140, c0_n6_w141, c0_n6_w142, c0_n6_w143, c0_n6_w144, c0_n6_w145, c0_n6_w146, c0_n6_w147, c0_n6_w148, c0_n6_w149, c0_n6_w150, c0_n6_w151, c0_n6_w152, c0_n6_w153, c0_n6_w154, c0_n6_w155, c0_n6_w156, c0_n6_w157, c0_n6_w158, c0_n6_w159, c0_n6_w160, c0_n6_w161, c0_n6_w162, c0_n6_w163, c0_n6_w164, c0_n6_w165, c0_n6_w166, c0_n6_w167, c0_n6_w168, c0_n6_w169, c0_n6_w170, c0_n6_w171, c0_n6_w172, c0_n6_w173, c0_n6_w174, c0_n6_w175, c0_n6_w176, c0_n6_w177, c0_n6_w178, c0_n6_w179, c0_n6_w180, c0_n6_w181, c0_n6_w182, c0_n6_w183, c0_n6_w184, c0_n6_w185, c0_n6_w186, c0_n6_w187, c0_n6_w188, c0_n6_w189, c0_n6_w190, c0_n6_w191, c0_n6_w192, c0_n6_w193, c0_n6_w194, c0_n6_w195, c0_n6_w196, c0_n6_w197, c0_n6_w198, c0_n6_w199, c0_n6_w200, c0_n7_w1, c0_n7_w2, c0_n7_w3, c0_n7_w4, c0_n7_w5, c0_n7_w6, c0_n7_w7, c0_n7_w8, c0_n7_w9, c0_n7_w10, c0_n7_w11, c0_n7_w12, c0_n7_w13, c0_n7_w14, c0_n7_w15, c0_n7_w16, c0_n7_w17, c0_n7_w18, c0_n7_w19, c0_n7_w20, c0_n7_w21, c0_n7_w22, c0_n7_w23, c0_n7_w24, c0_n7_w25, c0_n7_w26, c0_n7_w27, c0_n7_w28, c0_n7_w29, c0_n7_w30, c0_n7_w31, c0_n7_w32, c0_n7_w33, c0_n7_w34, c0_n7_w35, c0_n7_w36, c0_n7_w37, c0_n7_w38, c0_n7_w39, c0_n7_w40, c0_n7_w41, c0_n7_w42, c0_n7_w43, c0_n7_w44, c0_n7_w45, c0_n7_w46, c0_n7_w47, c0_n7_w48, c0_n7_w49, c0_n7_w50, c0_n7_w51, c0_n7_w52, c0_n7_w53, c0_n7_w54, c0_n7_w55, c0_n7_w56, c0_n7_w57, c0_n7_w58, c0_n7_w59, c0_n7_w60, c0_n7_w61, c0_n7_w62, c0_n7_w63, c0_n7_w64, c0_n7_w65, c0_n7_w66, c0_n7_w67, c0_n7_w68, c0_n7_w69, c0_n7_w70, c0_n7_w71, c0_n7_w72, c0_n7_w73, c0_n7_w74, c0_n7_w75, c0_n7_w76, c0_n7_w77, c0_n7_w78, c0_n7_w79, c0_n7_w80, c0_n7_w81, c0_n7_w82, c0_n7_w83, c0_n7_w84, c0_n7_w85, c0_n7_w86, c0_n7_w87, c0_n7_w88, c0_n7_w89, c0_n7_w90, c0_n7_w91, c0_n7_w92, c0_n7_w93, c0_n7_w94, c0_n7_w95, c0_n7_w96, c0_n7_w97, c0_n7_w98, c0_n7_w99, c0_n7_w100, c0_n7_w101, c0_n7_w102, c0_n7_w103, c0_n7_w104, c0_n7_w105, c0_n7_w106, c0_n7_w107, c0_n7_w108, c0_n7_w109, c0_n7_w110, c0_n7_w111, c0_n7_w112, c0_n7_w113, c0_n7_w114, c0_n7_w115, c0_n7_w116, c0_n7_w117, c0_n7_w118, c0_n7_w119, c0_n7_w120, c0_n7_w121, c0_n7_w122, c0_n7_w123, c0_n7_w124, c0_n7_w125, c0_n7_w126, c0_n7_w127, c0_n7_w128, c0_n7_w129, c0_n7_w130, c0_n7_w131, c0_n7_w132, c0_n7_w133, c0_n7_w134, c0_n7_w135, c0_n7_w136, c0_n7_w137, c0_n7_w138, c0_n7_w139, c0_n7_w140, c0_n7_w141, c0_n7_w142, c0_n7_w143, c0_n7_w144, c0_n7_w145, c0_n7_w146, c0_n7_w147, c0_n7_w148, c0_n7_w149, c0_n7_w150, c0_n7_w151, c0_n7_w152, c0_n7_w153, c0_n7_w154, c0_n7_w155, c0_n7_w156, c0_n7_w157, c0_n7_w158, c0_n7_w159, c0_n7_w160, c0_n7_w161, c0_n7_w162, c0_n7_w163, c0_n7_w164, c0_n7_w165, c0_n7_w166, c0_n7_w167, c0_n7_w168, c0_n7_w169, c0_n7_w170, c0_n7_w171, c0_n7_w172, c0_n7_w173, c0_n7_w174, c0_n7_w175, c0_n7_w176, c0_n7_w177, c0_n7_w178, c0_n7_w179, c0_n7_w180, c0_n7_w181, c0_n7_w182, c0_n7_w183, c0_n7_w184, c0_n7_w185, c0_n7_w186, c0_n7_w187, c0_n7_w188, c0_n7_w189, c0_n7_w190, c0_n7_w191, c0_n7_w192, c0_n7_w193, c0_n7_w194, c0_n7_w195, c0_n7_w196, c0_n7_w197, c0_n7_w198, c0_n7_w199, c0_n7_w200, c0_n8_w1, c0_n8_w2, c0_n8_w3, c0_n8_w4, c0_n8_w5, c0_n8_w6, c0_n8_w7, c0_n8_w8, c0_n8_w9, c0_n8_w10, c0_n8_w11, c0_n8_w12, c0_n8_w13, c0_n8_w14, c0_n8_w15, c0_n8_w16, c0_n8_w17, c0_n8_w18, c0_n8_w19, c0_n8_w20, c0_n8_w21, c0_n8_w22, c0_n8_w23, c0_n8_w24, c0_n8_w25, c0_n8_w26, c0_n8_w27, c0_n8_w28, c0_n8_w29, c0_n8_w30, c0_n8_w31, c0_n8_w32, c0_n8_w33, c0_n8_w34, c0_n8_w35, c0_n8_w36, c0_n8_w37, c0_n8_w38, c0_n8_w39, c0_n8_w40, c0_n8_w41, c0_n8_w42, c0_n8_w43, c0_n8_w44, c0_n8_w45, c0_n8_w46, c0_n8_w47, c0_n8_w48, c0_n8_w49, c0_n8_w50, c0_n8_w51, c0_n8_w52, c0_n8_w53, c0_n8_w54, c0_n8_w55, c0_n8_w56, c0_n8_w57, c0_n8_w58, c0_n8_w59, c0_n8_w60, c0_n8_w61, c0_n8_w62, c0_n8_w63, c0_n8_w64, c0_n8_w65, c0_n8_w66, c0_n8_w67, c0_n8_w68, c0_n8_w69, c0_n8_w70, c0_n8_w71, c0_n8_w72, c0_n8_w73, c0_n8_w74, c0_n8_w75, c0_n8_w76, c0_n8_w77, c0_n8_w78, c0_n8_w79, c0_n8_w80, c0_n8_w81, c0_n8_w82, c0_n8_w83, c0_n8_w84, c0_n8_w85, c0_n8_w86, c0_n8_w87, c0_n8_w88, c0_n8_w89, c0_n8_w90, c0_n8_w91, c0_n8_w92, c0_n8_w93, c0_n8_w94, c0_n8_w95, c0_n8_w96, c0_n8_w97, c0_n8_w98, c0_n8_w99, c0_n8_w100, c0_n8_w101, c0_n8_w102, c0_n8_w103, c0_n8_w104, c0_n8_w105, c0_n8_w106, c0_n8_w107, c0_n8_w108, c0_n8_w109, c0_n8_w110, c0_n8_w111, c0_n8_w112, c0_n8_w113, c0_n8_w114, c0_n8_w115, c0_n8_w116, c0_n8_w117, c0_n8_w118, c0_n8_w119, c0_n8_w120, c0_n8_w121, c0_n8_w122, c0_n8_w123, c0_n8_w124, c0_n8_w125, c0_n8_w126, c0_n8_w127, c0_n8_w128, c0_n8_w129, c0_n8_w130, c0_n8_w131, c0_n8_w132, c0_n8_w133, c0_n8_w134, c0_n8_w135, c0_n8_w136, c0_n8_w137, c0_n8_w138, c0_n8_w139, c0_n8_w140, c0_n8_w141, c0_n8_w142, c0_n8_w143, c0_n8_w144, c0_n8_w145, c0_n8_w146, c0_n8_w147, c0_n8_w148, c0_n8_w149, c0_n8_w150, c0_n8_w151, c0_n8_w152, c0_n8_w153, c0_n8_w154, c0_n8_w155, c0_n8_w156, c0_n8_w157, c0_n8_w158, c0_n8_w159, c0_n8_w160, c0_n8_w161, c0_n8_w162, c0_n8_w163, c0_n8_w164, c0_n8_w165, c0_n8_w166, c0_n8_w167, c0_n8_w168, c0_n8_w169, c0_n8_w170, c0_n8_w171, c0_n8_w172, c0_n8_w173, c0_n8_w174, c0_n8_w175, c0_n8_w176, c0_n8_w177, c0_n8_w178, c0_n8_w179, c0_n8_w180, c0_n8_w181, c0_n8_w182, c0_n8_w183, c0_n8_w184, c0_n8_w185, c0_n8_w186, c0_n8_w187, c0_n8_w188, c0_n8_w189, c0_n8_w190, c0_n8_w191, c0_n8_w192, c0_n8_w193, c0_n8_w194, c0_n8_w195, c0_n8_w196, c0_n8_w197, c0_n8_w198, c0_n8_w199, c0_n8_w200, c0_n9_w1, c0_n9_w2, c0_n9_w3, c0_n9_w4, c0_n9_w5, c0_n9_w6, c0_n9_w7, c0_n9_w8, c0_n9_w9, c0_n9_w10, c0_n9_w11, c0_n9_w12, c0_n9_w13, c0_n9_w14, c0_n9_w15, c0_n9_w16, c0_n9_w17, c0_n9_w18, c0_n9_w19, c0_n9_w20, c0_n9_w21, c0_n9_w22, c0_n9_w23, c0_n9_w24, c0_n9_w25, c0_n9_w26, c0_n9_w27, c0_n9_w28, c0_n9_w29, c0_n9_w30, c0_n9_w31, c0_n9_w32, c0_n9_w33, c0_n9_w34, c0_n9_w35, c0_n9_w36, c0_n9_w37, c0_n9_w38, c0_n9_w39, c0_n9_w40, c0_n9_w41, c0_n9_w42, c0_n9_w43, c0_n9_w44, c0_n9_w45, c0_n9_w46, c0_n9_w47, c0_n9_w48, c0_n9_w49, c0_n9_w50, c0_n9_w51, c0_n9_w52, c0_n9_w53, c0_n9_w54, c0_n9_w55, c0_n9_w56, c0_n9_w57, c0_n9_w58, c0_n9_w59, c0_n9_w60, c0_n9_w61, c0_n9_w62, c0_n9_w63, c0_n9_w64, c0_n9_w65, c0_n9_w66, c0_n9_w67, c0_n9_w68, c0_n9_w69, c0_n9_w70, c0_n9_w71, c0_n9_w72, c0_n9_w73, c0_n9_w74, c0_n9_w75, c0_n9_w76, c0_n9_w77, c0_n9_w78, c0_n9_w79, c0_n9_w80, c0_n9_w81, c0_n9_w82, c0_n9_w83, c0_n9_w84, c0_n9_w85, c0_n9_w86, c0_n9_w87, c0_n9_w88, c0_n9_w89, c0_n9_w90, c0_n9_w91, c0_n9_w92, c0_n9_w93, c0_n9_w94, c0_n9_w95, c0_n9_w96, c0_n9_w97, c0_n9_w98, c0_n9_w99, c0_n9_w100, c0_n9_w101, c0_n9_w102, c0_n9_w103, c0_n9_w104, c0_n9_w105, c0_n9_w106, c0_n9_w107, c0_n9_w108, c0_n9_w109, c0_n9_w110, c0_n9_w111, c0_n9_w112, c0_n9_w113, c0_n9_w114, c0_n9_w115, c0_n9_w116, c0_n9_w117, c0_n9_w118, c0_n9_w119, c0_n9_w120, c0_n9_w121, c0_n9_w122, c0_n9_w123, c0_n9_w124, c0_n9_w125, c0_n9_w126, c0_n9_w127, c0_n9_w128, c0_n9_w129, c0_n9_w130, c0_n9_w131, c0_n9_w132, c0_n9_w133, c0_n9_w134, c0_n9_w135, c0_n9_w136, c0_n9_w137, c0_n9_w138, c0_n9_w139, c0_n9_w140, c0_n9_w141, c0_n9_w142, c0_n9_w143, c0_n9_w144, c0_n9_w145, c0_n9_w146, c0_n9_w147, c0_n9_w148, c0_n9_w149, c0_n9_w150, c0_n9_w151, c0_n9_w152, c0_n9_w153, c0_n9_w154, c0_n9_w155, c0_n9_w156, c0_n9_w157, c0_n9_w158, c0_n9_w159, c0_n9_w160, c0_n9_w161, c0_n9_w162, c0_n9_w163, c0_n9_w164, c0_n9_w165, c0_n9_w166, c0_n9_w167, c0_n9_w168, c0_n9_w169, c0_n9_w170, c0_n9_w171, c0_n9_w172, c0_n9_w173, c0_n9_w174, c0_n9_w175, c0_n9_w176, c0_n9_w177, c0_n9_w178, c0_n9_w179, c0_n9_w180, c0_n9_w181, c0_n9_w182, c0_n9_w183, c0_n9_w184, c0_n9_w185, c0_n9_w186, c0_n9_w187, c0_n9_w188, c0_n9_w189, c0_n9_w190, c0_n9_w191, c0_n9_w192, c0_n9_w193, c0_n9_w194, c0_n9_w195, c0_n9_w196, c0_n9_w197, c0_n9_w198, c0_n9_w199, c0_n9_w200: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c0_n0_y, c0_n1_y, c0_n2_y, c0_n3_y, c0_n4_y, c0_n5_y, c0_n6_y, c0_n7_y, c0_n8_y, c0_n9_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada0_ReLU_10neuron_8bits_200n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n0_w1, 
            w2=> c0_n0_w2, 
            w3=> c0_n0_w3, 
            w4=> c0_n0_w4, 
            w5=> c0_n0_w5, 
            w6=> c0_n0_w6, 
            w7=> c0_n0_w7, 
            w8=> c0_n0_w8, 
            w9=> c0_n0_w9, 
            w10=> c0_n0_w10, 
            w11=> c0_n0_w11, 
            w12=> c0_n0_w12, 
            w13=> c0_n0_w13, 
            w14=> c0_n0_w14, 
            w15=> c0_n0_w15, 
            w16=> c0_n0_w16, 
            w17=> c0_n0_w17, 
            w18=> c0_n0_w18, 
            w19=> c0_n0_w19, 
            w20=> c0_n0_w20, 
            w21=> c0_n0_w21, 
            w22=> c0_n0_w22, 
            w23=> c0_n0_w23, 
            w24=> c0_n0_w24, 
            w25=> c0_n0_w25, 
            w26=> c0_n0_w26, 
            w27=> c0_n0_w27, 
            w28=> c0_n0_w28, 
            w29=> c0_n0_w29, 
            w30=> c0_n0_w30, 
            w31=> c0_n0_w31, 
            w32=> c0_n0_w32, 
            w33=> c0_n0_w33, 
            w34=> c0_n0_w34, 
            w35=> c0_n0_w35, 
            w36=> c0_n0_w36, 
            w37=> c0_n0_w37, 
            w38=> c0_n0_w38, 
            w39=> c0_n0_w39, 
            w40=> c0_n0_w40, 
            w41=> c0_n0_w41, 
            w42=> c0_n0_w42, 
            w43=> c0_n0_w43, 
            w44=> c0_n0_w44, 
            w45=> c0_n0_w45, 
            w46=> c0_n0_w46, 
            w47=> c0_n0_w47, 
            w48=> c0_n0_w48, 
            w49=> c0_n0_w49, 
            w50=> c0_n0_w50, 
            w51=> c0_n0_w51, 
            w52=> c0_n0_w52, 
            w53=> c0_n0_w53, 
            w54=> c0_n0_w54, 
            w55=> c0_n0_w55, 
            w56=> c0_n0_w56, 
            w57=> c0_n0_w57, 
            w58=> c0_n0_w58, 
            w59=> c0_n0_w59, 
            w60=> c0_n0_w60, 
            w61=> c0_n0_w61, 
            w62=> c0_n0_w62, 
            w63=> c0_n0_w63, 
            w64=> c0_n0_w64, 
            w65=> c0_n0_w65, 
            w66=> c0_n0_w66, 
            w67=> c0_n0_w67, 
            w68=> c0_n0_w68, 
            w69=> c0_n0_w69, 
            w70=> c0_n0_w70, 
            w71=> c0_n0_w71, 
            w72=> c0_n0_w72, 
            w73=> c0_n0_w73, 
            w74=> c0_n0_w74, 
            w75=> c0_n0_w75, 
            w76=> c0_n0_w76, 
            w77=> c0_n0_w77, 
            w78=> c0_n0_w78, 
            w79=> c0_n0_w79, 
            w80=> c0_n0_w80, 
            w81=> c0_n0_w81, 
            w82=> c0_n0_w82, 
            w83=> c0_n0_w83, 
            w84=> c0_n0_w84, 
            w85=> c0_n0_w85, 
            w86=> c0_n0_w86, 
            w87=> c0_n0_w87, 
            w88=> c0_n0_w88, 
            w89=> c0_n0_w89, 
            w90=> c0_n0_w90, 
            w91=> c0_n0_w91, 
            w92=> c0_n0_w92, 
            w93=> c0_n0_w93, 
            w94=> c0_n0_w94, 
            w95=> c0_n0_w95, 
            w96=> c0_n0_w96, 
            w97=> c0_n0_w97, 
            w98=> c0_n0_w98, 
            w99=> c0_n0_w99, 
            w100=> c0_n0_w100, 
            w101=> c0_n0_w101, 
            w102=> c0_n0_w102, 
            w103=> c0_n0_w103, 
            w104=> c0_n0_w104, 
            w105=> c0_n0_w105, 
            w106=> c0_n0_w106, 
            w107=> c0_n0_w107, 
            w108=> c0_n0_w108, 
            w109=> c0_n0_w109, 
            w110=> c0_n0_w110, 
            w111=> c0_n0_w111, 
            w112=> c0_n0_w112, 
            w113=> c0_n0_w113, 
            w114=> c0_n0_w114, 
            w115=> c0_n0_w115, 
            w116=> c0_n0_w116, 
            w117=> c0_n0_w117, 
            w118=> c0_n0_w118, 
            w119=> c0_n0_w119, 
            w120=> c0_n0_w120, 
            w121=> c0_n0_w121, 
            w122=> c0_n0_w122, 
            w123=> c0_n0_w123, 
            w124=> c0_n0_w124, 
            w125=> c0_n0_w125, 
            w126=> c0_n0_w126, 
            w127=> c0_n0_w127, 
            w128=> c0_n0_w128, 
            w129=> c0_n0_w129, 
            w130=> c0_n0_w130, 
            w131=> c0_n0_w131, 
            w132=> c0_n0_w132, 
            w133=> c0_n0_w133, 
            w134=> c0_n0_w134, 
            w135=> c0_n0_w135, 
            w136=> c0_n0_w136, 
            w137=> c0_n0_w137, 
            w138=> c0_n0_w138, 
            w139=> c0_n0_w139, 
            w140=> c0_n0_w140, 
            w141=> c0_n0_w141, 
            w142=> c0_n0_w142, 
            w143=> c0_n0_w143, 
            w144=> c0_n0_w144, 
            w145=> c0_n0_w145, 
            w146=> c0_n0_w146, 
            w147=> c0_n0_w147, 
            w148=> c0_n0_w148, 
            w149=> c0_n0_w149, 
            w150=> c0_n0_w150, 
            w151=> c0_n0_w151, 
            w152=> c0_n0_w152, 
            w153=> c0_n0_w153, 
            w154=> c0_n0_w154, 
            w155=> c0_n0_w155, 
            w156=> c0_n0_w156, 
            w157=> c0_n0_w157, 
            w158=> c0_n0_w158, 
            w159=> c0_n0_w159, 
            w160=> c0_n0_w160, 
            w161=> c0_n0_w161, 
            w162=> c0_n0_w162, 
            w163=> c0_n0_w163, 
            w164=> c0_n0_w164, 
            w165=> c0_n0_w165, 
            w166=> c0_n0_w166, 
            w167=> c0_n0_w167, 
            w168=> c0_n0_w168, 
            w169=> c0_n0_w169, 
            w170=> c0_n0_w170, 
            w171=> c0_n0_w171, 
            w172=> c0_n0_w172, 
            w173=> c0_n0_w173, 
            w174=> c0_n0_w174, 
            w175=> c0_n0_w175, 
            w176=> c0_n0_w176, 
            w177=> c0_n0_w177, 
            w178=> c0_n0_w178, 
            w179=> c0_n0_w179, 
            w180=> c0_n0_w180, 
            w181=> c0_n0_w181, 
            w182=> c0_n0_w182, 
            w183=> c0_n0_w183, 
            w184=> c0_n0_w184, 
            w185=> c0_n0_w185, 
            w186=> c0_n0_w186, 
            w187=> c0_n0_w187, 
            w188=> c0_n0_w188, 
            w189=> c0_n0_w189, 
            w190=> c0_n0_w190, 
            w191=> c0_n0_w191, 
            w192=> c0_n0_w192, 
            w193=> c0_n0_w193, 
            w194=> c0_n0_w194, 
            w195=> c0_n0_w195, 
            w196=> c0_n0_w196, 
            w197=> c0_n0_w197, 
            w198=> c0_n0_w198, 
            w199=> c0_n0_w199, 
            w200=> c0_n0_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n1_w1, 
            w2=> c0_n1_w2, 
            w3=> c0_n1_w3, 
            w4=> c0_n1_w4, 
            w5=> c0_n1_w5, 
            w6=> c0_n1_w6, 
            w7=> c0_n1_w7, 
            w8=> c0_n1_w8, 
            w9=> c0_n1_w9, 
            w10=> c0_n1_w10, 
            w11=> c0_n1_w11, 
            w12=> c0_n1_w12, 
            w13=> c0_n1_w13, 
            w14=> c0_n1_w14, 
            w15=> c0_n1_w15, 
            w16=> c0_n1_w16, 
            w17=> c0_n1_w17, 
            w18=> c0_n1_w18, 
            w19=> c0_n1_w19, 
            w20=> c0_n1_w20, 
            w21=> c0_n1_w21, 
            w22=> c0_n1_w22, 
            w23=> c0_n1_w23, 
            w24=> c0_n1_w24, 
            w25=> c0_n1_w25, 
            w26=> c0_n1_w26, 
            w27=> c0_n1_w27, 
            w28=> c0_n1_w28, 
            w29=> c0_n1_w29, 
            w30=> c0_n1_w30, 
            w31=> c0_n1_w31, 
            w32=> c0_n1_w32, 
            w33=> c0_n1_w33, 
            w34=> c0_n1_w34, 
            w35=> c0_n1_w35, 
            w36=> c0_n1_w36, 
            w37=> c0_n1_w37, 
            w38=> c0_n1_w38, 
            w39=> c0_n1_w39, 
            w40=> c0_n1_w40, 
            w41=> c0_n1_w41, 
            w42=> c0_n1_w42, 
            w43=> c0_n1_w43, 
            w44=> c0_n1_w44, 
            w45=> c0_n1_w45, 
            w46=> c0_n1_w46, 
            w47=> c0_n1_w47, 
            w48=> c0_n1_w48, 
            w49=> c0_n1_w49, 
            w50=> c0_n1_w50, 
            w51=> c0_n1_w51, 
            w52=> c0_n1_w52, 
            w53=> c0_n1_w53, 
            w54=> c0_n1_w54, 
            w55=> c0_n1_w55, 
            w56=> c0_n1_w56, 
            w57=> c0_n1_w57, 
            w58=> c0_n1_w58, 
            w59=> c0_n1_w59, 
            w60=> c0_n1_w60, 
            w61=> c0_n1_w61, 
            w62=> c0_n1_w62, 
            w63=> c0_n1_w63, 
            w64=> c0_n1_w64, 
            w65=> c0_n1_w65, 
            w66=> c0_n1_w66, 
            w67=> c0_n1_w67, 
            w68=> c0_n1_w68, 
            w69=> c0_n1_w69, 
            w70=> c0_n1_w70, 
            w71=> c0_n1_w71, 
            w72=> c0_n1_w72, 
            w73=> c0_n1_w73, 
            w74=> c0_n1_w74, 
            w75=> c0_n1_w75, 
            w76=> c0_n1_w76, 
            w77=> c0_n1_w77, 
            w78=> c0_n1_w78, 
            w79=> c0_n1_w79, 
            w80=> c0_n1_w80, 
            w81=> c0_n1_w81, 
            w82=> c0_n1_w82, 
            w83=> c0_n1_w83, 
            w84=> c0_n1_w84, 
            w85=> c0_n1_w85, 
            w86=> c0_n1_w86, 
            w87=> c0_n1_w87, 
            w88=> c0_n1_w88, 
            w89=> c0_n1_w89, 
            w90=> c0_n1_w90, 
            w91=> c0_n1_w91, 
            w92=> c0_n1_w92, 
            w93=> c0_n1_w93, 
            w94=> c0_n1_w94, 
            w95=> c0_n1_w95, 
            w96=> c0_n1_w96, 
            w97=> c0_n1_w97, 
            w98=> c0_n1_w98, 
            w99=> c0_n1_w99, 
            w100=> c0_n1_w100, 
            w101=> c0_n1_w101, 
            w102=> c0_n1_w102, 
            w103=> c0_n1_w103, 
            w104=> c0_n1_w104, 
            w105=> c0_n1_w105, 
            w106=> c0_n1_w106, 
            w107=> c0_n1_w107, 
            w108=> c0_n1_w108, 
            w109=> c0_n1_w109, 
            w110=> c0_n1_w110, 
            w111=> c0_n1_w111, 
            w112=> c0_n1_w112, 
            w113=> c0_n1_w113, 
            w114=> c0_n1_w114, 
            w115=> c0_n1_w115, 
            w116=> c0_n1_w116, 
            w117=> c0_n1_w117, 
            w118=> c0_n1_w118, 
            w119=> c0_n1_w119, 
            w120=> c0_n1_w120, 
            w121=> c0_n1_w121, 
            w122=> c0_n1_w122, 
            w123=> c0_n1_w123, 
            w124=> c0_n1_w124, 
            w125=> c0_n1_w125, 
            w126=> c0_n1_w126, 
            w127=> c0_n1_w127, 
            w128=> c0_n1_w128, 
            w129=> c0_n1_w129, 
            w130=> c0_n1_w130, 
            w131=> c0_n1_w131, 
            w132=> c0_n1_w132, 
            w133=> c0_n1_w133, 
            w134=> c0_n1_w134, 
            w135=> c0_n1_w135, 
            w136=> c0_n1_w136, 
            w137=> c0_n1_w137, 
            w138=> c0_n1_w138, 
            w139=> c0_n1_w139, 
            w140=> c0_n1_w140, 
            w141=> c0_n1_w141, 
            w142=> c0_n1_w142, 
            w143=> c0_n1_w143, 
            w144=> c0_n1_w144, 
            w145=> c0_n1_w145, 
            w146=> c0_n1_w146, 
            w147=> c0_n1_w147, 
            w148=> c0_n1_w148, 
            w149=> c0_n1_w149, 
            w150=> c0_n1_w150, 
            w151=> c0_n1_w151, 
            w152=> c0_n1_w152, 
            w153=> c0_n1_w153, 
            w154=> c0_n1_w154, 
            w155=> c0_n1_w155, 
            w156=> c0_n1_w156, 
            w157=> c0_n1_w157, 
            w158=> c0_n1_w158, 
            w159=> c0_n1_w159, 
            w160=> c0_n1_w160, 
            w161=> c0_n1_w161, 
            w162=> c0_n1_w162, 
            w163=> c0_n1_w163, 
            w164=> c0_n1_w164, 
            w165=> c0_n1_w165, 
            w166=> c0_n1_w166, 
            w167=> c0_n1_w167, 
            w168=> c0_n1_w168, 
            w169=> c0_n1_w169, 
            w170=> c0_n1_w170, 
            w171=> c0_n1_w171, 
            w172=> c0_n1_w172, 
            w173=> c0_n1_w173, 
            w174=> c0_n1_w174, 
            w175=> c0_n1_w175, 
            w176=> c0_n1_w176, 
            w177=> c0_n1_w177, 
            w178=> c0_n1_w178, 
            w179=> c0_n1_w179, 
            w180=> c0_n1_w180, 
            w181=> c0_n1_w181, 
            w182=> c0_n1_w182, 
            w183=> c0_n1_w183, 
            w184=> c0_n1_w184, 
            w185=> c0_n1_w185, 
            w186=> c0_n1_w186, 
            w187=> c0_n1_w187, 
            w188=> c0_n1_w188, 
            w189=> c0_n1_w189, 
            w190=> c0_n1_w190, 
            w191=> c0_n1_w191, 
            w192=> c0_n1_w192, 
            w193=> c0_n1_w193, 
            w194=> c0_n1_w194, 
            w195=> c0_n1_w195, 
            w196=> c0_n1_w196, 
            w197=> c0_n1_w197, 
            w198=> c0_n1_w198, 
            w199=> c0_n1_w199, 
            w200=> c0_n1_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n2_w1, 
            w2=> c0_n2_w2, 
            w3=> c0_n2_w3, 
            w4=> c0_n2_w4, 
            w5=> c0_n2_w5, 
            w6=> c0_n2_w6, 
            w7=> c0_n2_w7, 
            w8=> c0_n2_w8, 
            w9=> c0_n2_w9, 
            w10=> c0_n2_w10, 
            w11=> c0_n2_w11, 
            w12=> c0_n2_w12, 
            w13=> c0_n2_w13, 
            w14=> c0_n2_w14, 
            w15=> c0_n2_w15, 
            w16=> c0_n2_w16, 
            w17=> c0_n2_w17, 
            w18=> c0_n2_w18, 
            w19=> c0_n2_w19, 
            w20=> c0_n2_w20, 
            w21=> c0_n2_w21, 
            w22=> c0_n2_w22, 
            w23=> c0_n2_w23, 
            w24=> c0_n2_w24, 
            w25=> c0_n2_w25, 
            w26=> c0_n2_w26, 
            w27=> c0_n2_w27, 
            w28=> c0_n2_w28, 
            w29=> c0_n2_w29, 
            w30=> c0_n2_w30, 
            w31=> c0_n2_w31, 
            w32=> c0_n2_w32, 
            w33=> c0_n2_w33, 
            w34=> c0_n2_w34, 
            w35=> c0_n2_w35, 
            w36=> c0_n2_w36, 
            w37=> c0_n2_w37, 
            w38=> c0_n2_w38, 
            w39=> c0_n2_w39, 
            w40=> c0_n2_w40, 
            w41=> c0_n2_w41, 
            w42=> c0_n2_w42, 
            w43=> c0_n2_w43, 
            w44=> c0_n2_w44, 
            w45=> c0_n2_w45, 
            w46=> c0_n2_w46, 
            w47=> c0_n2_w47, 
            w48=> c0_n2_w48, 
            w49=> c0_n2_w49, 
            w50=> c0_n2_w50, 
            w51=> c0_n2_w51, 
            w52=> c0_n2_w52, 
            w53=> c0_n2_w53, 
            w54=> c0_n2_w54, 
            w55=> c0_n2_w55, 
            w56=> c0_n2_w56, 
            w57=> c0_n2_w57, 
            w58=> c0_n2_w58, 
            w59=> c0_n2_w59, 
            w60=> c0_n2_w60, 
            w61=> c0_n2_w61, 
            w62=> c0_n2_w62, 
            w63=> c0_n2_w63, 
            w64=> c0_n2_w64, 
            w65=> c0_n2_w65, 
            w66=> c0_n2_w66, 
            w67=> c0_n2_w67, 
            w68=> c0_n2_w68, 
            w69=> c0_n2_w69, 
            w70=> c0_n2_w70, 
            w71=> c0_n2_w71, 
            w72=> c0_n2_w72, 
            w73=> c0_n2_w73, 
            w74=> c0_n2_w74, 
            w75=> c0_n2_w75, 
            w76=> c0_n2_w76, 
            w77=> c0_n2_w77, 
            w78=> c0_n2_w78, 
            w79=> c0_n2_w79, 
            w80=> c0_n2_w80, 
            w81=> c0_n2_w81, 
            w82=> c0_n2_w82, 
            w83=> c0_n2_w83, 
            w84=> c0_n2_w84, 
            w85=> c0_n2_w85, 
            w86=> c0_n2_w86, 
            w87=> c0_n2_w87, 
            w88=> c0_n2_w88, 
            w89=> c0_n2_w89, 
            w90=> c0_n2_w90, 
            w91=> c0_n2_w91, 
            w92=> c0_n2_w92, 
            w93=> c0_n2_w93, 
            w94=> c0_n2_w94, 
            w95=> c0_n2_w95, 
            w96=> c0_n2_w96, 
            w97=> c0_n2_w97, 
            w98=> c0_n2_w98, 
            w99=> c0_n2_w99, 
            w100=> c0_n2_w100, 
            w101=> c0_n2_w101, 
            w102=> c0_n2_w102, 
            w103=> c0_n2_w103, 
            w104=> c0_n2_w104, 
            w105=> c0_n2_w105, 
            w106=> c0_n2_w106, 
            w107=> c0_n2_w107, 
            w108=> c0_n2_w108, 
            w109=> c0_n2_w109, 
            w110=> c0_n2_w110, 
            w111=> c0_n2_w111, 
            w112=> c0_n2_w112, 
            w113=> c0_n2_w113, 
            w114=> c0_n2_w114, 
            w115=> c0_n2_w115, 
            w116=> c0_n2_w116, 
            w117=> c0_n2_w117, 
            w118=> c0_n2_w118, 
            w119=> c0_n2_w119, 
            w120=> c0_n2_w120, 
            w121=> c0_n2_w121, 
            w122=> c0_n2_w122, 
            w123=> c0_n2_w123, 
            w124=> c0_n2_w124, 
            w125=> c0_n2_w125, 
            w126=> c0_n2_w126, 
            w127=> c0_n2_w127, 
            w128=> c0_n2_w128, 
            w129=> c0_n2_w129, 
            w130=> c0_n2_w130, 
            w131=> c0_n2_w131, 
            w132=> c0_n2_w132, 
            w133=> c0_n2_w133, 
            w134=> c0_n2_w134, 
            w135=> c0_n2_w135, 
            w136=> c0_n2_w136, 
            w137=> c0_n2_w137, 
            w138=> c0_n2_w138, 
            w139=> c0_n2_w139, 
            w140=> c0_n2_w140, 
            w141=> c0_n2_w141, 
            w142=> c0_n2_w142, 
            w143=> c0_n2_w143, 
            w144=> c0_n2_w144, 
            w145=> c0_n2_w145, 
            w146=> c0_n2_w146, 
            w147=> c0_n2_w147, 
            w148=> c0_n2_w148, 
            w149=> c0_n2_w149, 
            w150=> c0_n2_w150, 
            w151=> c0_n2_w151, 
            w152=> c0_n2_w152, 
            w153=> c0_n2_w153, 
            w154=> c0_n2_w154, 
            w155=> c0_n2_w155, 
            w156=> c0_n2_w156, 
            w157=> c0_n2_w157, 
            w158=> c0_n2_w158, 
            w159=> c0_n2_w159, 
            w160=> c0_n2_w160, 
            w161=> c0_n2_w161, 
            w162=> c0_n2_w162, 
            w163=> c0_n2_w163, 
            w164=> c0_n2_w164, 
            w165=> c0_n2_w165, 
            w166=> c0_n2_w166, 
            w167=> c0_n2_w167, 
            w168=> c0_n2_w168, 
            w169=> c0_n2_w169, 
            w170=> c0_n2_w170, 
            w171=> c0_n2_w171, 
            w172=> c0_n2_w172, 
            w173=> c0_n2_w173, 
            w174=> c0_n2_w174, 
            w175=> c0_n2_w175, 
            w176=> c0_n2_w176, 
            w177=> c0_n2_w177, 
            w178=> c0_n2_w178, 
            w179=> c0_n2_w179, 
            w180=> c0_n2_w180, 
            w181=> c0_n2_w181, 
            w182=> c0_n2_w182, 
            w183=> c0_n2_w183, 
            w184=> c0_n2_w184, 
            w185=> c0_n2_w185, 
            w186=> c0_n2_w186, 
            w187=> c0_n2_w187, 
            w188=> c0_n2_w188, 
            w189=> c0_n2_w189, 
            w190=> c0_n2_w190, 
            w191=> c0_n2_w191, 
            w192=> c0_n2_w192, 
            w193=> c0_n2_w193, 
            w194=> c0_n2_w194, 
            w195=> c0_n2_w195, 
            w196=> c0_n2_w196, 
            w197=> c0_n2_w197, 
            w198=> c0_n2_w198, 
            w199=> c0_n2_w199, 
            w200=> c0_n2_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n3_w1, 
            w2=> c0_n3_w2, 
            w3=> c0_n3_w3, 
            w4=> c0_n3_w4, 
            w5=> c0_n3_w5, 
            w6=> c0_n3_w6, 
            w7=> c0_n3_w7, 
            w8=> c0_n3_w8, 
            w9=> c0_n3_w9, 
            w10=> c0_n3_w10, 
            w11=> c0_n3_w11, 
            w12=> c0_n3_w12, 
            w13=> c0_n3_w13, 
            w14=> c0_n3_w14, 
            w15=> c0_n3_w15, 
            w16=> c0_n3_w16, 
            w17=> c0_n3_w17, 
            w18=> c0_n3_w18, 
            w19=> c0_n3_w19, 
            w20=> c0_n3_w20, 
            w21=> c0_n3_w21, 
            w22=> c0_n3_w22, 
            w23=> c0_n3_w23, 
            w24=> c0_n3_w24, 
            w25=> c0_n3_w25, 
            w26=> c0_n3_w26, 
            w27=> c0_n3_w27, 
            w28=> c0_n3_w28, 
            w29=> c0_n3_w29, 
            w30=> c0_n3_w30, 
            w31=> c0_n3_w31, 
            w32=> c0_n3_w32, 
            w33=> c0_n3_w33, 
            w34=> c0_n3_w34, 
            w35=> c0_n3_w35, 
            w36=> c0_n3_w36, 
            w37=> c0_n3_w37, 
            w38=> c0_n3_w38, 
            w39=> c0_n3_w39, 
            w40=> c0_n3_w40, 
            w41=> c0_n3_w41, 
            w42=> c0_n3_w42, 
            w43=> c0_n3_w43, 
            w44=> c0_n3_w44, 
            w45=> c0_n3_w45, 
            w46=> c0_n3_w46, 
            w47=> c0_n3_w47, 
            w48=> c0_n3_w48, 
            w49=> c0_n3_w49, 
            w50=> c0_n3_w50, 
            w51=> c0_n3_w51, 
            w52=> c0_n3_w52, 
            w53=> c0_n3_w53, 
            w54=> c0_n3_w54, 
            w55=> c0_n3_w55, 
            w56=> c0_n3_w56, 
            w57=> c0_n3_w57, 
            w58=> c0_n3_w58, 
            w59=> c0_n3_w59, 
            w60=> c0_n3_w60, 
            w61=> c0_n3_w61, 
            w62=> c0_n3_w62, 
            w63=> c0_n3_w63, 
            w64=> c0_n3_w64, 
            w65=> c0_n3_w65, 
            w66=> c0_n3_w66, 
            w67=> c0_n3_w67, 
            w68=> c0_n3_w68, 
            w69=> c0_n3_w69, 
            w70=> c0_n3_w70, 
            w71=> c0_n3_w71, 
            w72=> c0_n3_w72, 
            w73=> c0_n3_w73, 
            w74=> c0_n3_w74, 
            w75=> c0_n3_w75, 
            w76=> c0_n3_w76, 
            w77=> c0_n3_w77, 
            w78=> c0_n3_w78, 
            w79=> c0_n3_w79, 
            w80=> c0_n3_w80, 
            w81=> c0_n3_w81, 
            w82=> c0_n3_w82, 
            w83=> c0_n3_w83, 
            w84=> c0_n3_w84, 
            w85=> c0_n3_w85, 
            w86=> c0_n3_w86, 
            w87=> c0_n3_w87, 
            w88=> c0_n3_w88, 
            w89=> c0_n3_w89, 
            w90=> c0_n3_w90, 
            w91=> c0_n3_w91, 
            w92=> c0_n3_w92, 
            w93=> c0_n3_w93, 
            w94=> c0_n3_w94, 
            w95=> c0_n3_w95, 
            w96=> c0_n3_w96, 
            w97=> c0_n3_w97, 
            w98=> c0_n3_w98, 
            w99=> c0_n3_w99, 
            w100=> c0_n3_w100, 
            w101=> c0_n3_w101, 
            w102=> c0_n3_w102, 
            w103=> c0_n3_w103, 
            w104=> c0_n3_w104, 
            w105=> c0_n3_w105, 
            w106=> c0_n3_w106, 
            w107=> c0_n3_w107, 
            w108=> c0_n3_w108, 
            w109=> c0_n3_w109, 
            w110=> c0_n3_w110, 
            w111=> c0_n3_w111, 
            w112=> c0_n3_w112, 
            w113=> c0_n3_w113, 
            w114=> c0_n3_w114, 
            w115=> c0_n3_w115, 
            w116=> c0_n3_w116, 
            w117=> c0_n3_w117, 
            w118=> c0_n3_w118, 
            w119=> c0_n3_w119, 
            w120=> c0_n3_w120, 
            w121=> c0_n3_w121, 
            w122=> c0_n3_w122, 
            w123=> c0_n3_w123, 
            w124=> c0_n3_w124, 
            w125=> c0_n3_w125, 
            w126=> c0_n3_w126, 
            w127=> c0_n3_w127, 
            w128=> c0_n3_w128, 
            w129=> c0_n3_w129, 
            w130=> c0_n3_w130, 
            w131=> c0_n3_w131, 
            w132=> c0_n3_w132, 
            w133=> c0_n3_w133, 
            w134=> c0_n3_w134, 
            w135=> c0_n3_w135, 
            w136=> c0_n3_w136, 
            w137=> c0_n3_w137, 
            w138=> c0_n3_w138, 
            w139=> c0_n3_w139, 
            w140=> c0_n3_w140, 
            w141=> c0_n3_w141, 
            w142=> c0_n3_w142, 
            w143=> c0_n3_w143, 
            w144=> c0_n3_w144, 
            w145=> c0_n3_w145, 
            w146=> c0_n3_w146, 
            w147=> c0_n3_w147, 
            w148=> c0_n3_w148, 
            w149=> c0_n3_w149, 
            w150=> c0_n3_w150, 
            w151=> c0_n3_w151, 
            w152=> c0_n3_w152, 
            w153=> c0_n3_w153, 
            w154=> c0_n3_w154, 
            w155=> c0_n3_w155, 
            w156=> c0_n3_w156, 
            w157=> c0_n3_w157, 
            w158=> c0_n3_w158, 
            w159=> c0_n3_w159, 
            w160=> c0_n3_w160, 
            w161=> c0_n3_w161, 
            w162=> c0_n3_w162, 
            w163=> c0_n3_w163, 
            w164=> c0_n3_w164, 
            w165=> c0_n3_w165, 
            w166=> c0_n3_w166, 
            w167=> c0_n3_w167, 
            w168=> c0_n3_w168, 
            w169=> c0_n3_w169, 
            w170=> c0_n3_w170, 
            w171=> c0_n3_w171, 
            w172=> c0_n3_w172, 
            w173=> c0_n3_w173, 
            w174=> c0_n3_w174, 
            w175=> c0_n3_w175, 
            w176=> c0_n3_w176, 
            w177=> c0_n3_w177, 
            w178=> c0_n3_w178, 
            w179=> c0_n3_w179, 
            w180=> c0_n3_w180, 
            w181=> c0_n3_w181, 
            w182=> c0_n3_w182, 
            w183=> c0_n3_w183, 
            w184=> c0_n3_w184, 
            w185=> c0_n3_w185, 
            w186=> c0_n3_w186, 
            w187=> c0_n3_w187, 
            w188=> c0_n3_w188, 
            w189=> c0_n3_w189, 
            w190=> c0_n3_w190, 
            w191=> c0_n3_w191, 
            w192=> c0_n3_w192, 
            w193=> c0_n3_w193, 
            w194=> c0_n3_w194, 
            w195=> c0_n3_w195, 
            w196=> c0_n3_w196, 
            w197=> c0_n3_w197, 
            w198=> c0_n3_w198, 
            w199=> c0_n3_w199, 
            w200=> c0_n3_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n4_w1, 
            w2=> c0_n4_w2, 
            w3=> c0_n4_w3, 
            w4=> c0_n4_w4, 
            w5=> c0_n4_w5, 
            w6=> c0_n4_w6, 
            w7=> c0_n4_w7, 
            w8=> c0_n4_w8, 
            w9=> c0_n4_w9, 
            w10=> c0_n4_w10, 
            w11=> c0_n4_w11, 
            w12=> c0_n4_w12, 
            w13=> c0_n4_w13, 
            w14=> c0_n4_w14, 
            w15=> c0_n4_w15, 
            w16=> c0_n4_w16, 
            w17=> c0_n4_w17, 
            w18=> c0_n4_w18, 
            w19=> c0_n4_w19, 
            w20=> c0_n4_w20, 
            w21=> c0_n4_w21, 
            w22=> c0_n4_w22, 
            w23=> c0_n4_w23, 
            w24=> c0_n4_w24, 
            w25=> c0_n4_w25, 
            w26=> c0_n4_w26, 
            w27=> c0_n4_w27, 
            w28=> c0_n4_w28, 
            w29=> c0_n4_w29, 
            w30=> c0_n4_w30, 
            w31=> c0_n4_w31, 
            w32=> c0_n4_w32, 
            w33=> c0_n4_w33, 
            w34=> c0_n4_w34, 
            w35=> c0_n4_w35, 
            w36=> c0_n4_w36, 
            w37=> c0_n4_w37, 
            w38=> c0_n4_w38, 
            w39=> c0_n4_w39, 
            w40=> c0_n4_w40, 
            w41=> c0_n4_w41, 
            w42=> c0_n4_w42, 
            w43=> c0_n4_w43, 
            w44=> c0_n4_w44, 
            w45=> c0_n4_w45, 
            w46=> c0_n4_w46, 
            w47=> c0_n4_w47, 
            w48=> c0_n4_w48, 
            w49=> c0_n4_w49, 
            w50=> c0_n4_w50, 
            w51=> c0_n4_w51, 
            w52=> c0_n4_w52, 
            w53=> c0_n4_w53, 
            w54=> c0_n4_w54, 
            w55=> c0_n4_w55, 
            w56=> c0_n4_w56, 
            w57=> c0_n4_w57, 
            w58=> c0_n4_w58, 
            w59=> c0_n4_w59, 
            w60=> c0_n4_w60, 
            w61=> c0_n4_w61, 
            w62=> c0_n4_w62, 
            w63=> c0_n4_w63, 
            w64=> c0_n4_w64, 
            w65=> c0_n4_w65, 
            w66=> c0_n4_w66, 
            w67=> c0_n4_w67, 
            w68=> c0_n4_w68, 
            w69=> c0_n4_w69, 
            w70=> c0_n4_w70, 
            w71=> c0_n4_w71, 
            w72=> c0_n4_w72, 
            w73=> c0_n4_w73, 
            w74=> c0_n4_w74, 
            w75=> c0_n4_w75, 
            w76=> c0_n4_w76, 
            w77=> c0_n4_w77, 
            w78=> c0_n4_w78, 
            w79=> c0_n4_w79, 
            w80=> c0_n4_w80, 
            w81=> c0_n4_w81, 
            w82=> c0_n4_w82, 
            w83=> c0_n4_w83, 
            w84=> c0_n4_w84, 
            w85=> c0_n4_w85, 
            w86=> c0_n4_w86, 
            w87=> c0_n4_w87, 
            w88=> c0_n4_w88, 
            w89=> c0_n4_w89, 
            w90=> c0_n4_w90, 
            w91=> c0_n4_w91, 
            w92=> c0_n4_w92, 
            w93=> c0_n4_w93, 
            w94=> c0_n4_w94, 
            w95=> c0_n4_w95, 
            w96=> c0_n4_w96, 
            w97=> c0_n4_w97, 
            w98=> c0_n4_w98, 
            w99=> c0_n4_w99, 
            w100=> c0_n4_w100, 
            w101=> c0_n4_w101, 
            w102=> c0_n4_w102, 
            w103=> c0_n4_w103, 
            w104=> c0_n4_w104, 
            w105=> c0_n4_w105, 
            w106=> c0_n4_w106, 
            w107=> c0_n4_w107, 
            w108=> c0_n4_w108, 
            w109=> c0_n4_w109, 
            w110=> c0_n4_w110, 
            w111=> c0_n4_w111, 
            w112=> c0_n4_w112, 
            w113=> c0_n4_w113, 
            w114=> c0_n4_w114, 
            w115=> c0_n4_w115, 
            w116=> c0_n4_w116, 
            w117=> c0_n4_w117, 
            w118=> c0_n4_w118, 
            w119=> c0_n4_w119, 
            w120=> c0_n4_w120, 
            w121=> c0_n4_w121, 
            w122=> c0_n4_w122, 
            w123=> c0_n4_w123, 
            w124=> c0_n4_w124, 
            w125=> c0_n4_w125, 
            w126=> c0_n4_w126, 
            w127=> c0_n4_w127, 
            w128=> c0_n4_w128, 
            w129=> c0_n4_w129, 
            w130=> c0_n4_w130, 
            w131=> c0_n4_w131, 
            w132=> c0_n4_w132, 
            w133=> c0_n4_w133, 
            w134=> c0_n4_w134, 
            w135=> c0_n4_w135, 
            w136=> c0_n4_w136, 
            w137=> c0_n4_w137, 
            w138=> c0_n4_w138, 
            w139=> c0_n4_w139, 
            w140=> c0_n4_w140, 
            w141=> c0_n4_w141, 
            w142=> c0_n4_w142, 
            w143=> c0_n4_w143, 
            w144=> c0_n4_w144, 
            w145=> c0_n4_w145, 
            w146=> c0_n4_w146, 
            w147=> c0_n4_w147, 
            w148=> c0_n4_w148, 
            w149=> c0_n4_w149, 
            w150=> c0_n4_w150, 
            w151=> c0_n4_w151, 
            w152=> c0_n4_w152, 
            w153=> c0_n4_w153, 
            w154=> c0_n4_w154, 
            w155=> c0_n4_w155, 
            w156=> c0_n4_w156, 
            w157=> c0_n4_w157, 
            w158=> c0_n4_w158, 
            w159=> c0_n4_w159, 
            w160=> c0_n4_w160, 
            w161=> c0_n4_w161, 
            w162=> c0_n4_w162, 
            w163=> c0_n4_w163, 
            w164=> c0_n4_w164, 
            w165=> c0_n4_w165, 
            w166=> c0_n4_w166, 
            w167=> c0_n4_w167, 
            w168=> c0_n4_w168, 
            w169=> c0_n4_w169, 
            w170=> c0_n4_w170, 
            w171=> c0_n4_w171, 
            w172=> c0_n4_w172, 
            w173=> c0_n4_w173, 
            w174=> c0_n4_w174, 
            w175=> c0_n4_w175, 
            w176=> c0_n4_w176, 
            w177=> c0_n4_w177, 
            w178=> c0_n4_w178, 
            w179=> c0_n4_w179, 
            w180=> c0_n4_w180, 
            w181=> c0_n4_w181, 
            w182=> c0_n4_w182, 
            w183=> c0_n4_w183, 
            w184=> c0_n4_w184, 
            w185=> c0_n4_w185, 
            w186=> c0_n4_w186, 
            w187=> c0_n4_w187, 
            w188=> c0_n4_w188, 
            w189=> c0_n4_w189, 
            w190=> c0_n4_w190, 
            w191=> c0_n4_w191, 
            w192=> c0_n4_w192, 
            w193=> c0_n4_w193, 
            w194=> c0_n4_w194, 
            w195=> c0_n4_w195, 
            w196=> c0_n4_w196, 
            w197=> c0_n4_w197, 
            w198=> c0_n4_w198, 
            w199=> c0_n4_w199, 
            w200=> c0_n4_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n5_w1, 
            w2=> c0_n5_w2, 
            w3=> c0_n5_w3, 
            w4=> c0_n5_w4, 
            w5=> c0_n5_w5, 
            w6=> c0_n5_w6, 
            w7=> c0_n5_w7, 
            w8=> c0_n5_w8, 
            w9=> c0_n5_w9, 
            w10=> c0_n5_w10, 
            w11=> c0_n5_w11, 
            w12=> c0_n5_w12, 
            w13=> c0_n5_w13, 
            w14=> c0_n5_w14, 
            w15=> c0_n5_w15, 
            w16=> c0_n5_w16, 
            w17=> c0_n5_w17, 
            w18=> c0_n5_w18, 
            w19=> c0_n5_w19, 
            w20=> c0_n5_w20, 
            w21=> c0_n5_w21, 
            w22=> c0_n5_w22, 
            w23=> c0_n5_w23, 
            w24=> c0_n5_w24, 
            w25=> c0_n5_w25, 
            w26=> c0_n5_w26, 
            w27=> c0_n5_w27, 
            w28=> c0_n5_w28, 
            w29=> c0_n5_w29, 
            w30=> c0_n5_w30, 
            w31=> c0_n5_w31, 
            w32=> c0_n5_w32, 
            w33=> c0_n5_w33, 
            w34=> c0_n5_w34, 
            w35=> c0_n5_w35, 
            w36=> c0_n5_w36, 
            w37=> c0_n5_w37, 
            w38=> c0_n5_w38, 
            w39=> c0_n5_w39, 
            w40=> c0_n5_w40, 
            w41=> c0_n5_w41, 
            w42=> c0_n5_w42, 
            w43=> c0_n5_w43, 
            w44=> c0_n5_w44, 
            w45=> c0_n5_w45, 
            w46=> c0_n5_w46, 
            w47=> c0_n5_w47, 
            w48=> c0_n5_w48, 
            w49=> c0_n5_w49, 
            w50=> c0_n5_w50, 
            w51=> c0_n5_w51, 
            w52=> c0_n5_w52, 
            w53=> c0_n5_w53, 
            w54=> c0_n5_w54, 
            w55=> c0_n5_w55, 
            w56=> c0_n5_w56, 
            w57=> c0_n5_w57, 
            w58=> c0_n5_w58, 
            w59=> c0_n5_w59, 
            w60=> c0_n5_w60, 
            w61=> c0_n5_w61, 
            w62=> c0_n5_w62, 
            w63=> c0_n5_w63, 
            w64=> c0_n5_w64, 
            w65=> c0_n5_w65, 
            w66=> c0_n5_w66, 
            w67=> c0_n5_w67, 
            w68=> c0_n5_w68, 
            w69=> c0_n5_w69, 
            w70=> c0_n5_w70, 
            w71=> c0_n5_w71, 
            w72=> c0_n5_w72, 
            w73=> c0_n5_w73, 
            w74=> c0_n5_w74, 
            w75=> c0_n5_w75, 
            w76=> c0_n5_w76, 
            w77=> c0_n5_w77, 
            w78=> c0_n5_w78, 
            w79=> c0_n5_w79, 
            w80=> c0_n5_w80, 
            w81=> c0_n5_w81, 
            w82=> c0_n5_w82, 
            w83=> c0_n5_w83, 
            w84=> c0_n5_w84, 
            w85=> c0_n5_w85, 
            w86=> c0_n5_w86, 
            w87=> c0_n5_w87, 
            w88=> c0_n5_w88, 
            w89=> c0_n5_w89, 
            w90=> c0_n5_w90, 
            w91=> c0_n5_w91, 
            w92=> c0_n5_w92, 
            w93=> c0_n5_w93, 
            w94=> c0_n5_w94, 
            w95=> c0_n5_w95, 
            w96=> c0_n5_w96, 
            w97=> c0_n5_w97, 
            w98=> c0_n5_w98, 
            w99=> c0_n5_w99, 
            w100=> c0_n5_w100, 
            w101=> c0_n5_w101, 
            w102=> c0_n5_w102, 
            w103=> c0_n5_w103, 
            w104=> c0_n5_w104, 
            w105=> c0_n5_w105, 
            w106=> c0_n5_w106, 
            w107=> c0_n5_w107, 
            w108=> c0_n5_w108, 
            w109=> c0_n5_w109, 
            w110=> c0_n5_w110, 
            w111=> c0_n5_w111, 
            w112=> c0_n5_w112, 
            w113=> c0_n5_w113, 
            w114=> c0_n5_w114, 
            w115=> c0_n5_w115, 
            w116=> c0_n5_w116, 
            w117=> c0_n5_w117, 
            w118=> c0_n5_w118, 
            w119=> c0_n5_w119, 
            w120=> c0_n5_w120, 
            w121=> c0_n5_w121, 
            w122=> c0_n5_w122, 
            w123=> c0_n5_w123, 
            w124=> c0_n5_w124, 
            w125=> c0_n5_w125, 
            w126=> c0_n5_w126, 
            w127=> c0_n5_w127, 
            w128=> c0_n5_w128, 
            w129=> c0_n5_w129, 
            w130=> c0_n5_w130, 
            w131=> c0_n5_w131, 
            w132=> c0_n5_w132, 
            w133=> c0_n5_w133, 
            w134=> c0_n5_w134, 
            w135=> c0_n5_w135, 
            w136=> c0_n5_w136, 
            w137=> c0_n5_w137, 
            w138=> c0_n5_w138, 
            w139=> c0_n5_w139, 
            w140=> c0_n5_w140, 
            w141=> c0_n5_w141, 
            w142=> c0_n5_w142, 
            w143=> c0_n5_w143, 
            w144=> c0_n5_w144, 
            w145=> c0_n5_w145, 
            w146=> c0_n5_w146, 
            w147=> c0_n5_w147, 
            w148=> c0_n5_w148, 
            w149=> c0_n5_w149, 
            w150=> c0_n5_w150, 
            w151=> c0_n5_w151, 
            w152=> c0_n5_w152, 
            w153=> c0_n5_w153, 
            w154=> c0_n5_w154, 
            w155=> c0_n5_w155, 
            w156=> c0_n5_w156, 
            w157=> c0_n5_w157, 
            w158=> c0_n5_w158, 
            w159=> c0_n5_w159, 
            w160=> c0_n5_w160, 
            w161=> c0_n5_w161, 
            w162=> c0_n5_w162, 
            w163=> c0_n5_w163, 
            w164=> c0_n5_w164, 
            w165=> c0_n5_w165, 
            w166=> c0_n5_w166, 
            w167=> c0_n5_w167, 
            w168=> c0_n5_w168, 
            w169=> c0_n5_w169, 
            w170=> c0_n5_w170, 
            w171=> c0_n5_w171, 
            w172=> c0_n5_w172, 
            w173=> c0_n5_w173, 
            w174=> c0_n5_w174, 
            w175=> c0_n5_w175, 
            w176=> c0_n5_w176, 
            w177=> c0_n5_w177, 
            w178=> c0_n5_w178, 
            w179=> c0_n5_w179, 
            w180=> c0_n5_w180, 
            w181=> c0_n5_w181, 
            w182=> c0_n5_w182, 
            w183=> c0_n5_w183, 
            w184=> c0_n5_w184, 
            w185=> c0_n5_w185, 
            w186=> c0_n5_w186, 
            w187=> c0_n5_w187, 
            w188=> c0_n5_w188, 
            w189=> c0_n5_w189, 
            w190=> c0_n5_w190, 
            w191=> c0_n5_w191, 
            w192=> c0_n5_w192, 
            w193=> c0_n5_w193, 
            w194=> c0_n5_w194, 
            w195=> c0_n5_w195, 
            w196=> c0_n5_w196, 
            w197=> c0_n5_w197, 
            w198=> c0_n5_w198, 
            w199=> c0_n5_w199, 
            w200=> c0_n5_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n6_w1, 
            w2=> c0_n6_w2, 
            w3=> c0_n6_w3, 
            w4=> c0_n6_w4, 
            w5=> c0_n6_w5, 
            w6=> c0_n6_w6, 
            w7=> c0_n6_w7, 
            w8=> c0_n6_w8, 
            w9=> c0_n6_w9, 
            w10=> c0_n6_w10, 
            w11=> c0_n6_w11, 
            w12=> c0_n6_w12, 
            w13=> c0_n6_w13, 
            w14=> c0_n6_w14, 
            w15=> c0_n6_w15, 
            w16=> c0_n6_w16, 
            w17=> c0_n6_w17, 
            w18=> c0_n6_w18, 
            w19=> c0_n6_w19, 
            w20=> c0_n6_w20, 
            w21=> c0_n6_w21, 
            w22=> c0_n6_w22, 
            w23=> c0_n6_w23, 
            w24=> c0_n6_w24, 
            w25=> c0_n6_w25, 
            w26=> c0_n6_w26, 
            w27=> c0_n6_w27, 
            w28=> c0_n6_w28, 
            w29=> c0_n6_w29, 
            w30=> c0_n6_w30, 
            w31=> c0_n6_w31, 
            w32=> c0_n6_w32, 
            w33=> c0_n6_w33, 
            w34=> c0_n6_w34, 
            w35=> c0_n6_w35, 
            w36=> c0_n6_w36, 
            w37=> c0_n6_w37, 
            w38=> c0_n6_w38, 
            w39=> c0_n6_w39, 
            w40=> c0_n6_w40, 
            w41=> c0_n6_w41, 
            w42=> c0_n6_w42, 
            w43=> c0_n6_w43, 
            w44=> c0_n6_w44, 
            w45=> c0_n6_w45, 
            w46=> c0_n6_w46, 
            w47=> c0_n6_w47, 
            w48=> c0_n6_w48, 
            w49=> c0_n6_w49, 
            w50=> c0_n6_w50, 
            w51=> c0_n6_w51, 
            w52=> c0_n6_w52, 
            w53=> c0_n6_w53, 
            w54=> c0_n6_w54, 
            w55=> c0_n6_w55, 
            w56=> c0_n6_w56, 
            w57=> c0_n6_w57, 
            w58=> c0_n6_w58, 
            w59=> c0_n6_w59, 
            w60=> c0_n6_w60, 
            w61=> c0_n6_w61, 
            w62=> c0_n6_w62, 
            w63=> c0_n6_w63, 
            w64=> c0_n6_w64, 
            w65=> c0_n6_w65, 
            w66=> c0_n6_w66, 
            w67=> c0_n6_w67, 
            w68=> c0_n6_w68, 
            w69=> c0_n6_w69, 
            w70=> c0_n6_w70, 
            w71=> c0_n6_w71, 
            w72=> c0_n6_w72, 
            w73=> c0_n6_w73, 
            w74=> c0_n6_w74, 
            w75=> c0_n6_w75, 
            w76=> c0_n6_w76, 
            w77=> c0_n6_w77, 
            w78=> c0_n6_w78, 
            w79=> c0_n6_w79, 
            w80=> c0_n6_w80, 
            w81=> c0_n6_w81, 
            w82=> c0_n6_w82, 
            w83=> c0_n6_w83, 
            w84=> c0_n6_w84, 
            w85=> c0_n6_w85, 
            w86=> c0_n6_w86, 
            w87=> c0_n6_w87, 
            w88=> c0_n6_w88, 
            w89=> c0_n6_w89, 
            w90=> c0_n6_w90, 
            w91=> c0_n6_w91, 
            w92=> c0_n6_w92, 
            w93=> c0_n6_w93, 
            w94=> c0_n6_w94, 
            w95=> c0_n6_w95, 
            w96=> c0_n6_w96, 
            w97=> c0_n6_w97, 
            w98=> c0_n6_w98, 
            w99=> c0_n6_w99, 
            w100=> c0_n6_w100, 
            w101=> c0_n6_w101, 
            w102=> c0_n6_w102, 
            w103=> c0_n6_w103, 
            w104=> c0_n6_w104, 
            w105=> c0_n6_w105, 
            w106=> c0_n6_w106, 
            w107=> c0_n6_w107, 
            w108=> c0_n6_w108, 
            w109=> c0_n6_w109, 
            w110=> c0_n6_w110, 
            w111=> c0_n6_w111, 
            w112=> c0_n6_w112, 
            w113=> c0_n6_w113, 
            w114=> c0_n6_w114, 
            w115=> c0_n6_w115, 
            w116=> c0_n6_w116, 
            w117=> c0_n6_w117, 
            w118=> c0_n6_w118, 
            w119=> c0_n6_w119, 
            w120=> c0_n6_w120, 
            w121=> c0_n6_w121, 
            w122=> c0_n6_w122, 
            w123=> c0_n6_w123, 
            w124=> c0_n6_w124, 
            w125=> c0_n6_w125, 
            w126=> c0_n6_w126, 
            w127=> c0_n6_w127, 
            w128=> c0_n6_w128, 
            w129=> c0_n6_w129, 
            w130=> c0_n6_w130, 
            w131=> c0_n6_w131, 
            w132=> c0_n6_w132, 
            w133=> c0_n6_w133, 
            w134=> c0_n6_w134, 
            w135=> c0_n6_w135, 
            w136=> c0_n6_w136, 
            w137=> c0_n6_w137, 
            w138=> c0_n6_w138, 
            w139=> c0_n6_w139, 
            w140=> c0_n6_w140, 
            w141=> c0_n6_w141, 
            w142=> c0_n6_w142, 
            w143=> c0_n6_w143, 
            w144=> c0_n6_w144, 
            w145=> c0_n6_w145, 
            w146=> c0_n6_w146, 
            w147=> c0_n6_w147, 
            w148=> c0_n6_w148, 
            w149=> c0_n6_w149, 
            w150=> c0_n6_w150, 
            w151=> c0_n6_w151, 
            w152=> c0_n6_w152, 
            w153=> c0_n6_w153, 
            w154=> c0_n6_w154, 
            w155=> c0_n6_w155, 
            w156=> c0_n6_w156, 
            w157=> c0_n6_w157, 
            w158=> c0_n6_w158, 
            w159=> c0_n6_w159, 
            w160=> c0_n6_w160, 
            w161=> c0_n6_w161, 
            w162=> c0_n6_w162, 
            w163=> c0_n6_w163, 
            w164=> c0_n6_w164, 
            w165=> c0_n6_w165, 
            w166=> c0_n6_w166, 
            w167=> c0_n6_w167, 
            w168=> c0_n6_w168, 
            w169=> c0_n6_w169, 
            w170=> c0_n6_w170, 
            w171=> c0_n6_w171, 
            w172=> c0_n6_w172, 
            w173=> c0_n6_w173, 
            w174=> c0_n6_w174, 
            w175=> c0_n6_w175, 
            w176=> c0_n6_w176, 
            w177=> c0_n6_w177, 
            w178=> c0_n6_w178, 
            w179=> c0_n6_w179, 
            w180=> c0_n6_w180, 
            w181=> c0_n6_w181, 
            w182=> c0_n6_w182, 
            w183=> c0_n6_w183, 
            w184=> c0_n6_w184, 
            w185=> c0_n6_w185, 
            w186=> c0_n6_w186, 
            w187=> c0_n6_w187, 
            w188=> c0_n6_w188, 
            w189=> c0_n6_w189, 
            w190=> c0_n6_w190, 
            w191=> c0_n6_w191, 
            w192=> c0_n6_w192, 
            w193=> c0_n6_w193, 
            w194=> c0_n6_w194, 
            w195=> c0_n6_w195, 
            w196=> c0_n6_w196, 
            w197=> c0_n6_w197, 
            w198=> c0_n6_w198, 
            w199=> c0_n6_w199, 
            w200=> c0_n6_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n7_w1, 
            w2=> c0_n7_w2, 
            w3=> c0_n7_w3, 
            w4=> c0_n7_w4, 
            w5=> c0_n7_w5, 
            w6=> c0_n7_w6, 
            w7=> c0_n7_w7, 
            w8=> c0_n7_w8, 
            w9=> c0_n7_w9, 
            w10=> c0_n7_w10, 
            w11=> c0_n7_w11, 
            w12=> c0_n7_w12, 
            w13=> c0_n7_w13, 
            w14=> c0_n7_w14, 
            w15=> c0_n7_w15, 
            w16=> c0_n7_w16, 
            w17=> c0_n7_w17, 
            w18=> c0_n7_w18, 
            w19=> c0_n7_w19, 
            w20=> c0_n7_w20, 
            w21=> c0_n7_w21, 
            w22=> c0_n7_w22, 
            w23=> c0_n7_w23, 
            w24=> c0_n7_w24, 
            w25=> c0_n7_w25, 
            w26=> c0_n7_w26, 
            w27=> c0_n7_w27, 
            w28=> c0_n7_w28, 
            w29=> c0_n7_w29, 
            w30=> c0_n7_w30, 
            w31=> c0_n7_w31, 
            w32=> c0_n7_w32, 
            w33=> c0_n7_w33, 
            w34=> c0_n7_w34, 
            w35=> c0_n7_w35, 
            w36=> c0_n7_w36, 
            w37=> c0_n7_w37, 
            w38=> c0_n7_w38, 
            w39=> c0_n7_w39, 
            w40=> c0_n7_w40, 
            w41=> c0_n7_w41, 
            w42=> c0_n7_w42, 
            w43=> c0_n7_w43, 
            w44=> c0_n7_w44, 
            w45=> c0_n7_w45, 
            w46=> c0_n7_w46, 
            w47=> c0_n7_w47, 
            w48=> c0_n7_w48, 
            w49=> c0_n7_w49, 
            w50=> c0_n7_w50, 
            w51=> c0_n7_w51, 
            w52=> c0_n7_w52, 
            w53=> c0_n7_w53, 
            w54=> c0_n7_w54, 
            w55=> c0_n7_w55, 
            w56=> c0_n7_w56, 
            w57=> c0_n7_w57, 
            w58=> c0_n7_w58, 
            w59=> c0_n7_w59, 
            w60=> c0_n7_w60, 
            w61=> c0_n7_w61, 
            w62=> c0_n7_w62, 
            w63=> c0_n7_w63, 
            w64=> c0_n7_w64, 
            w65=> c0_n7_w65, 
            w66=> c0_n7_w66, 
            w67=> c0_n7_w67, 
            w68=> c0_n7_w68, 
            w69=> c0_n7_w69, 
            w70=> c0_n7_w70, 
            w71=> c0_n7_w71, 
            w72=> c0_n7_w72, 
            w73=> c0_n7_w73, 
            w74=> c0_n7_w74, 
            w75=> c0_n7_w75, 
            w76=> c0_n7_w76, 
            w77=> c0_n7_w77, 
            w78=> c0_n7_w78, 
            w79=> c0_n7_w79, 
            w80=> c0_n7_w80, 
            w81=> c0_n7_w81, 
            w82=> c0_n7_w82, 
            w83=> c0_n7_w83, 
            w84=> c0_n7_w84, 
            w85=> c0_n7_w85, 
            w86=> c0_n7_w86, 
            w87=> c0_n7_w87, 
            w88=> c0_n7_w88, 
            w89=> c0_n7_w89, 
            w90=> c0_n7_w90, 
            w91=> c0_n7_w91, 
            w92=> c0_n7_w92, 
            w93=> c0_n7_w93, 
            w94=> c0_n7_w94, 
            w95=> c0_n7_w95, 
            w96=> c0_n7_w96, 
            w97=> c0_n7_w97, 
            w98=> c0_n7_w98, 
            w99=> c0_n7_w99, 
            w100=> c0_n7_w100, 
            w101=> c0_n7_w101, 
            w102=> c0_n7_w102, 
            w103=> c0_n7_w103, 
            w104=> c0_n7_w104, 
            w105=> c0_n7_w105, 
            w106=> c0_n7_w106, 
            w107=> c0_n7_w107, 
            w108=> c0_n7_w108, 
            w109=> c0_n7_w109, 
            w110=> c0_n7_w110, 
            w111=> c0_n7_w111, 
            w112=> c0_n7_w112, 
            w113=> c0_n7_w113, 
            w114=> c0_n7_w114, 
            w115=> c0_n7_w115, 
            w116=> c0_n7_w116, 
            w117=> c0_n7_w117, 
            w118=> c0_n7_w118, 
            w119=> c0_n7_w119, 
            w120=> c0_n7_w120, 
            w121=> c0_n7_w121, 
            w122=> c0_n7_w122, 
            w123=> c0_n7_w123, 
            w124=> c0_n7_w124, 
            w125=> c0_n7_w125, 
            w126=> c0_n7_w126, 
            w127=> c0_n7_w127, 
            w128=> c0_n7_w128, 
            w129=> c0_n7_w129, 
            w130=> c0_n7_w130, 
            w131=> c0_n7_w131, 
            w132=> c0_n7_w132, 
            w133=> c0_n7_w133, 
            w134=> c0_n7_w134, 
            w135=> c0_n7_w135, 
            w136=> c0_n7_w136, 
            w137=> c0_n7_w137, 
            w138=> c0_n7_w138, 
            w139=> c0_n7_w139, 
            w140=> c0_n7_w140, 
            w141=> c0_n7_w141, 
            w142=> c0_n7_w142, 
            w143=> c0_n7_w143, 
            w144=> c0_n7_w144, 
            w145=> c0_n7_w145, 
            w146=> c0_n7_w146, 
            w147=> c0_n7_w147, 
            w148=> c0_n7_w148, 
            w149=> c0_n7_w149, 
            w150=> c0_n7_w150, 
            w151=> c0_n7_w151, 
            w152=> c0_n7_w152, 
            w153=> c0_n7_w153, 
            w154=> c0_n7_w154, 
            w155=> c0_n7_w155, 
            w156=> c0_n7_w156, 
            w157=> c0_n7_w157, 
            w158=> c0_n7_w158, 
            w159=> c0_n7_w159, 
            w160=> c0_n7_w160, 
            w161=> c0_n7_w161, 
            w162=> c0_n7_w162, 
            w163=> c0_n7_w163, 
            w164=> c0_n7_w164, 
            w165=> c0_n7_w165, 
            w166=> c0_n7_w166, 
            w167=> c0_n7_w167, 
            w168=> c0_n7_w168, 
            w169=> c0_n7_w169, 
            w170=> c0_n7_w170, 
            w171=> c0_n7_w171, 
            w172=> c0_n7_w172, 
            w173=> c0_n7_w173, 
            w174=> c0_n7_w174, 
            w175=> c0_n7_w175, 
            w176=> c0_n7_w176, 
            w177=> c0_n7_w177, 
            w178=> c0_n7_w178, 
            w179=> c0_n7_w179, 
            w180=> c0_n7_w180, 
            w181=> c0_n7_w181, 
            w182=> c0_n7_w182, 
            w183=> c0_n7_w183, 
            w184=> c0_n7_w184, 
            w185=> c0_n7_w185, 
            w186=> c0_n7_w186, 
            w187=> c0_n7_w187, 
            w188=> c0_n7_w188, 
            w189=> c0_n7_w189, 
            w190=> c0_n7_w190, 
            w191=> c0_n7_w191, 
            w192=> c0_n7_w192, 
            w193=> c0_n7_w193, 
            w194=> c0_n7_w194, 
            w195=> c0_n7_w195, 
            w196=> c0_n7_w196, 
            w197=> c0_n7_w197, 
            w198=> c0_n7_w198, 
            w199=> c0_n7_w199, 
            w200=> c0_n7_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n8_w1, 
            w2=> c0_n8_w2, 
            w3=> c0_n8_w3, 
            w4=> c0_n8_w4, 
            w5=> c0_n8_w5, 
            w6=> c0_n8_w6, 
            w7=> c0_n8_w7, 
            w8=> c0_n8_w8, 
            w9=> c0_n8_w9, 
            w10=> c0_n8_w10, 
            w11=> c0_n8_w11, 
            w12=> c0_n8_w12, 
            w13=> c0_n8_w13, 
            w14=> c0_n8_w14, 
            w15=> c0_n8_w15, 
            w16=> c0_n8_w16, 
            w17=> c0_n8_w17, 
            w18=> c0_n8_w18, 
            w19=> c0_n8_w19, 
            w20=> c0_n8_w20, 
            w21=> c0_n8_w21, 
            w22=> c0_n8_w22, 
            w23=> c0_n8_w23, 
            w24=> c0_n8_w24, 
            w25=> c0_n8_w25, 
            w26=> c0_n8_w26, 
            w27=> c0_n8_w27, 
            w28=> c0_n8_w28, 
            w29=> c0_n8_w29, 
            w30=> c0_n8_w30, 
            w31=> c0_n8_w31, 
            w32=> c0_n8_w32, 
            w33=> c0_n8_w33, 
            w34=> c0_n8_w34, 
            w35=> c0_n8_w35, 
            w36=> c0_n8_w36, 
            w37=> c0_n8_w37, 
            w38=> c0_n8_w38, 
            w39=> c0_n8_w39, 
            w40=> c0_n8_w40, 
            w41=> c0_n8_w41, 
            w42=> c0_n8_w42, 
            w43=> c0_n8_w43, 
            w44=> c0_n8_w44, 
            w45=> c0_n8_w45, 
            w46=> c0_n8_w46, 
            w47=> c0_n8_w47, 
            w48=> c0_n8_w48, 
            w49=> c0_n8_w49, 
            w50=> c0_n8_w50, 
            w51=> c0_n8_w51, 
            w52=> c0_n8_w52, 
            w53=> c0_n8_w53, 
            w54=> c0_n8_w54, 
            w55=> c0_n8_w55, 
            w56=> c0_n8_w56, 
            w57=> c0_n8_w57, 
            w58=> c0_n8_w58, 
            w59=> c0_n8_w59, 
            w60=> c0_n8_w60, 
            w61=> c0_n8_w61, 
            w62=> c0_n8_w62, 
            w63=> c0_n8_w63, 
            w64=> c0_n8_w64, 
            w65=> c0_n8_w65, 
            w66=> c0_n8_w66, 
            w67=> c0_n8_w67, 
            w68=> c0_n8_w68, 
            w69=> c0_n8_w69, 
            w70=> c0_n8_w70, 
            w71=> c0_n8_w71, 
            w72=> c0_n8_w72, 
            w73=> c0_n8_w73, 
            w74=> c0_n8_w74, 
            w75=> c0_n8_w75, 
            w76=> c0_n8_w76, 
            w77=> c0_n8_w77, 
            w78=> c0_n8_w78, 
            w79=> c0_n8_w79, 
            w80=> c0_n8_w80, 
            w81=> c0_n8_w81, 
            w82=> c0_n8_w82, 
            w83=> c0_n8_w83, 
            w84=> c0_n8_w84, 
            w85=> c0_n8_w85, 
            w86=> c0_n8_w86, 
            w87=> c0_n8_w87, 
            w88=> c0_n8_w88, 
            w89=> c0_n8_w89, 
            w90=> c0_n8_w90, 
            w91=> c0_n8_w91, 
            w92=> c0_n8_w92, 
            w93=> c0_n8_w93, 
            w94=> c0_n8_w94, 
            w95=> c0_n8_w95, 
            w96=> c0_n8_w96, 
            w97=> c0_n8_w97, 
            w98=> c0_n8_w98, 
            w99=> c0_n8_w99, 
            w100=> c0_n8_w100, 
            w101=> c0_n8_w101, 
            w102=> c0_n8_w102, 
            w103=> c0_n8_w103, 
            w104=> c0_n8_w104, 
            w105=> c0_n8_w105, 
            w106=> c0_n8_w106, 
            w107=> c0_n8_w107, 
            w108=> c0_n8_w108, 
            w109=> c0_n8_w109, 
            w110=> c0_n8_w110, 
            w111=> c0_n8_w111, 
            w112=> c0_n8_w112, 
            w113=> c0_n8_w113, 
            w114=> c0_n8_w114, 
            w115=> c0_n8_w115, 
            w116=> c0_n8_w116, 
            w117=> c0_n8_w117, 
            w118=> c0_n8_w118, 
            w119=> c0_n8_w119, 
            w120=> c0_n8_w120, 
            w121=> c0_n8_w121, 
            w122=> c0_n8_w122, 
            w123=> c0_n8_w123, 
            w124=> c0_n8_w124, 
            w125=> c0_n8_w125, 
            w126=> c0_n8_w126, 
            w127=> c0_n8_w127, 
            w128=> c0_n8_w128, 
            w129=> c0_n8_w129, 
            w130=> c0_n8_w130, 
            w131=> c0_n8_w131, 
            w132=> c0_n8_w132, 
            w133=> c0_n8_w133, 
            w134=> c0_n8_w134, 
            w135=> c0_n8_w135, 
            w136=> c0_n8_w136, 
            w137=> c0_n8_w137, 
            w138=> c0_n8_w138, 
            w139=> c0_n8_w139, 
            w140=> c0_n8_w140, 
            w141=> c0_n8_w141, 
            w142=> c0_n8_w142, 
            w143=> c0_n8_w143, 
            w144=> c0_n8_w144, 
            w145=> c0_n8_w145, 
            w146=> c0_n8_w146, 
            w147=> c0_n8_w147, 
            w148=> c0_n8_w148, 
            w149=> c0_n8_w149, 
            w150=> c0_n8_w150, 
            w151=> c0_n8_w151, 
            w152=> c0_n8_w152, 
            w153=> c0_n8_w153, 
            w154=> c0_n8_w154, 
            w155=> c0_n8_w155, 
            w156=> c0_n8_w156, 
            w157=> c0_n8_w157, 
            w158=> c0_n8_w158, 
            w159=> c0_n8_w159, 
            w160=> c0_n8_w160, 
            w161=> c0_n8_w161, 
            w162=> c0_n8_w162, 
            w163=> c0_n8_w163, 
            w164=> c0_n8_w164, 
            w165=> c0_n8_w165, 
            w166=> c0_n8_w166, 
            w167=> c0_n8_w167, 
            w168=> c0_n8_w168, 
            w169=> c0_n8_w169, 
            w170=> c0_n8_w170, 
            w171=> c0_n8_w171, 
            w172=> c0_n8_w172, 
            w173=> c0_n8_w173, 
            w174=> c0_n8_w174, 
            w175=> c0_n8_w175, 
            w176=> c0_n8_w176, 
            w177=> c0_n8_w177, 
            w178=> c0_n8_w178, 
            w179=> c0_n8_w179, 
            w180=> c0_n8_w180, 
            w181=> c0_n8_w181, 
            w182=> c0_n8_w182, 
            w183=> c0_n8_w183, 
            w184=> c0_n8_w184, 
            w185=> c0_n8_w185, 
            w186=> c0_n8_w186, 
            w187=> c0_n8_w187, 
            w188=> c0_n8_w188, 
            w189=> c0_n8_w189, 
            w190=> c0_n8_w190, 
            w191=> c0_n8_w191, 
            w192=> c0_n8_w192, 
            w193=> c0_n8_w193, 
            w194=> c0_n8_w194, 
            w195=> c0_n8_w195, 
            w196=> c0_n8_w196, 
            w197=> c0_n8_w197, 
            w198=> c0_n8_w198, 
            w199=> c0_n8_w199, 
            w200=> c0_n8_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_ReLU_200n_8bit_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n9_w1, 
            w2=> c0_n9_w2, 
            w3=> c0_n9_w3, 
            w4=> c0_n9_w4, 
            w5=> c0_n9_w5, 
            w6=> c0_n9_w6, 
            w7=> c0_n9_w7, 
            w8=> c0_n9_w8, 
            w9=> c0_n9_w9, 
            w10=> c0_n9_w10, 
            w11=> c0_n9_w11, 
            w12=> c0_n9_w12, 
            w13=> c0_n9_w13, 
            w14=> c0_n9_w14, 
            w15=> c0_n9_w15, 
            w16=> c0_n9_w16, 
            w17=> c0_n9_w17, 
            w18=> c0_n9_w18, 
            w19=> c0_n9_w19, 
            w20=> c0_n9_w20, 
            w21=> c0_n9_w21, 
            w22=> c0_n9_w22, 
            w23=> c0_n9_w23, 
            w24=> c0_n9_w24, 
            w25=> c0_n9_w25, 
            w26=> c0_n9_w26, 
            w27=> c0_n9_w27, 
            w28=> c0_n9_w28, 
            w29=> c0_n9_w29, 
            w30=> c0_n9_w30, 
            w31=> c0_n9_w31, 
            w32=> c0_n9_w32, 
            w33=> c0_n9_w33, 
            w34=> c0_n9_w34, 
            w35=> c0_n9_w35, 
            w36=> c0_n9_w36, 
            w37=> c0_n9_w37, 
            w38=> c0_n9_w38, 
            w39=> c0_n9_w39, 
            w40=> c0_n9_w40, 
            w41=> c0_n9_w41, 
            w42=> c0_n9_w42, 
            w43=> c0_n9_w43, 
            w44=> c0_n9_w44, 
            w45=> c0_n9_w45, 
            w46=> c0_n9_w46, 
            w47=> c0_n9_w47, 
            w48=> c0_n9_w48, 
            w49=> c0_n9_w49, 
            w50=> c0_n9_w50, 
            w51=> c0_n9_w51, 
            w52=> c0_n9_w52, 
            w53=> c0_n9_w53, 
            w54=> c0_n9_w54, 
            w55=> c0_n9_w55, 
            w56=> c0_n9_w56, 
            w57=> c0_n9_w57, 
            w58=> c0_n9_w58, 
            w59=> c0_n9_w59, 
            w60=> c0_n9_w60, 
            w61=> c0_n9_w61, 
            w62=> c0_n9_w62, 
            w63=> c0_n9_w63, 
            w64=> c0_n9_w64, 
            w65=> c0_n9_w65, 
            w66=> c0_n9_w66, 
            w67=> c0_n9_w67, 
            w68=> c0_n9_w68, 
            w69=> c0_n9_w69, 
            w70=> c0_n9_w70, 
            w71=> c0_n9_w71, 
            w72=> c0_n9_w72, 
            w73=> c0_n9_w73, 
            w74=> c0_n9_w74, 
            w75=> c0_n9_w75, 
            w76=> c0_n9_w76, 
            w77=> c0_n9_w77, 
            w78=> c0_n9_w78, 
            w79=> c0_n9_w79, 
            w80=> c0_n9_w80, 
            w81=> c0_n9_w81, 
            w82=> c0_n9_w82, 
            w83=> c0_n9_w83, 
            w84=> c0_n9_w84, 
            w85=> c0_n9_w85, 
            w86=> c0_n9_w86, 
            w87=> c0_n9_w87, 
            w88=> c0_n9_w88, 
            w89=> c0_n9_w89, 
            w90=> c0_n9_w90, 
            w91=> c0_n9_w91, 
            w92=> c0_n9_w92, 
            w93=> c0_n9_w93, 
            w94=> c0_n9_w94, 
            w95=> c0_n9_w95, 
            w96=> c0_n9_w96, 
            w97=> c0_n9_w97, 
            w98=> c0_n9_w98, 
            w99=> c0_n9_w99, 
            w100=> c0_n9_w100, 
            w101=> c0_n9_w101, 
            w102=> c0_n9_w102, 
            w103=> c0_n9_w103, 
            w104=> c0_n9_w104, 
            w105=> c0_n9_w105, 
            w106=> c0_n9_w106, 
            w107=> c0_n9_w107, 
            w108=> c0_n9_w108, 
            w109=> c0_n9_w109, 
            w110=> c0_n9_w110, 
            w111=> c0_n9_w111, 
            w112=> c0_n9_w112, 
            w113=> c0_n9_w113, 
            w114=> c0_n9_w114, 
            w115=> c0_n9_w115, 
            w116=> c0_n9_w116, 
            w117=> c0_n9_w117, 
            w118=> c0_n9_w118, 
            w119=> c0_n9_w119, 
            w120=> c0_n9_w120, 
            w121=> c0_n9_w121, 
            w122=> c0_n9_w122, 
            w123=> c0_n9_w123, 
            w124=> c0_n9_w124, 
            w125=> c0_n9_w125, 
            w126=> c0_n9_w126, 
            w127=> c0_n9_w127, 
            w128=> c0_n9_w128, 
            w129=> c0_n9_w129, 
            w130=> c0_n9_w130, 
            w131=> c0_n9_w131, 
            w132=> c0_n9_w132, 
            w133=> c0_n9_w133, 
            w134=> c0_n9_w134, 
            w135=> c0_n9_w135, 
            w136=> c0_n9_w136, 
            w137=> c0_n9_w137, 
            w138=> c0_n9_w138, 
            w139=> c0_n9_w139, 
            w140=> c0_n9_w140, 
            w141=> c0_n9_w141, 
            w142=> c0_n9_w142, 
            w143=> c0_n9_w143, 
            w144=> c0_n9_w144, 
            w145=> c0_n9_w145, 
            w146=> c0_n9_w146, 
            w147=> c0_n9_w147, 
            w148=> c0_n9_w148, 
            w149=> c0_n9_w149, 
            w150=> c0_n9_w150, 
            w151=> c0_n9_w151, 
            w152=> c0_n9_w152, 
            w153=> c0_n9_w153, 
            w154=> c0_n9_w154, 
            w155=> c0_n9_w155, 
            w156=> c0_n9_w156, 
            w157=> c0_n9_w157, 
            w158=> c0_n9_w158, 
            w159=> c0_n9_w159, 
            w160=> c0_n9_w160, 
            w161=> c0_n9_w161, 
            w162=> c0_n9_w162, 
            w163=> c0_n9_w163, 
            w164=> c0_n9_w164, 
            w165=> c0_n9_w165, 
            w166=> c0_n9_w166, 
            w167=> c0_n9_w167, 
            w168=> c0_n9_w168, 
            w169=> c0_n9_w169, 
            w170=> c0_n9_w170, 
            w171=> c0_n9_w171, 
            w172=> c0_n9_w172, 
            w173=> c0_n9_w173, 
            w174=> c0_n9_w174, 
            w175=> c0_n9_w175, 
            w176=> c0_n9_w176, 
            w177=> c0_n9_w177, 
            w178=> c0_n9_w178, 
            w179=> c0_n9_w179, 
            w180=> c0_n9_w180, 
            w181=> c0_n9_w181, 
            w182=> c0_n9_w182, 
            w183=> c0_n9_w183, 
            w184=> c0_n9_w184, 
            w185=> c0_n9_w185, 
            w186=> c0_n9_w186, 
            w187=> c0_n9_w187, 
            w188=> c0_n9_w188, 
            w189=> c0_n9_w189, 
            w190=> c0_n9_w190, 
            w191=> c0_n9_w191, 
            w192=> c0_n9_w192, 
            w193=> c0_n9_w193, 
            w194=> c0_n9_w194, 
            w195=> c0_n9_w195, 
            w196=> c0_n9_w196, 
            w197=> c0_n9_w197, 
            w198=> c0_n9_w198, 
            w199=> c0_n9_w199, 
            w200=> c0_n9_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n9_y
   );           
             
END ARCHITECTURE;
