LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada0_ReLU_100neuron_8bits_200n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c0_n0_bias, c0_n1_bias, c0_n2_bias, c0_n3_bias, c0_n4_bias, c0_n5_bias, c0_n6_bias, c0_n7_bias, c0_n8_bias, c0_n9_bias, c0_n10_bias, c0_n11_bias, c0_n12_bias, c0_n13_bias, c0_n14_bias, c0_n15_bias, c0_n16_bias, c0_n17_bias, c0_n18_bias, c0_n19_bias, c0_n20_bias, c0_n21_bias, c0_n22_bias, c0_n23_bias, c0_n24_bias, c0_n25_bias, c0_n26_bias, c0_n27_bias, c0_n28_bias, c0_n29_bias, c0_n30_bias, c0_n31_bias, c0_n32_bias, c0_n33_bias, c0_n34_bias, c0_n35_bias, c0_n36_bias, c0_n37_bias, c0_n38_bias, c0_n39_bias, c0_n40_bias, c0_n41_bias, c0_n42_bias, c0_n43_bias, c0_n44_bias, c0_n45_bias, c0_n46_bias, c0_n47_bias, c0_n48_bias, c0_n49_bias, c0_n50_bias, c0_n51_bias, c0_n52_bias, c0_n53_bias, c0_n54_bias, c0_n55_bias, c0_n56_bias, c0_n57_bias, c0_n58_bias, c0_n59_bias, c0_n60_bias, c0_n61_bias, c0_n62_bias, c0_n63_bias, c0_n64_bias, c0_n65_bias, c0_n66_bias, c0_n67_bias, c0_n68_bias, c0_n69_bias, c0_n70_bias, c0_n71_bias, c0_n72_bias, c0_n73_bias, c0_n74_bias, c0_n75_bias, c0_n76_bias, c0_n77_bias, c0_n78_bias, c0_n79_bias, c0_n80_bias, c0_n81_bias, c0_n82_bias, c0_n83_bias, c0_n84_bias, c0_n85_bias, c0_n86_bias, c0_n87_bias, c0_n88_bias, c0_n89_bias, c0_n90_bias, c0_n91_bias, c0_n92_bias, c0_n93_bias, c0_n94_bias, c0_n95_bias, c0_n96_bias, c0_n97_bias, c0_n98_bias, c0_n99_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, c0_n0_w1, c0_n0_w2, c0_n0_w3, c0_n0_w4, c0_n0_w5, c0_n0_w6, c0_n0_w7, c0_n0_w8, c0_n0_w9, c0_n0_w10, c0_n0_w11, c0_n0_w12, c0_n0_w13, c0_n0_w14, c0_n0_w15, c0_n0_w16, c0_n0_w17, c0_n0_w18, c0_n0_w19, c0_n0_w20, c0_n0_w21, c0_n0_w22, c0_n0_w23, c0_n0_w24, c0_n0_w25, c0_n0_w26, c0_n0_w27, c0_n0_w28, c0_n0_w29, c0_n0_w30, c0_n0_w31, c0_n0_w32, c0_n0_w33, c0_n0_w34, c0_n0_w35, c0_n0_w36, c0_n0_w37, c0_n0_w38, c0_n0_w39, c0_n0_w40, c0_n0_w41, c0_n0_w42, c0_n0_w43, c0_n0_w44, c0_n0_w45, c0_n0_w46, c0_n0_w47, c0_n0_w48, c0_n0_w49, c0_n0_w50, c0_n0_w51, c0_n0_w52, c0_n0_w53, c0_n0_w54, c0_n0_w55, c0_n0_w56, c0_n0_w57, c0_n0_w58, c0_n0_w59, c0_n0_w60, c0_n0_w61, c0_n0_w62, c0_n0_w63, c0_n0_w64, c0_n0_w65, c0_n0_w66, c0_n0_w67, c0_n0_w68, c0_n0_w69, c0_n0_w70, c0_n0_w71, c0_n0_w72, c0_n0_w73, c0_n0_w74, c0_n0_w75, c0_n0_w76, c0_n0_w77, c0_n0_w78, c0_n0_w79, c0_n0_w80, c0_n0_w81, c0_n0_w82, c0_n0_w83, c0_n0_w84, c0_n0_w85, c0_n0_w86, c0_n0_w87, c0_n0_w88, c0_n0_w89, c0_n0_w90, c0_n0_w91, c0_n0_w92, c0_n0_w93, c0_n0_w94, c0_n0_w95, c0_n0_w96, c0_n0_w97, c0_n0_w98, c0_n0_w99, c0_n0_w100, c0_n0_w101, c0_n0_w102, c0_n0_w103, c0_n0_w104, c0_n0_w105, c0_n0_w106, c0_n0_w107, c0_n0_w108, c0_n0_w109, c0_n0_w110, c0_n0_w111, c0_n0_w112, c0_n0_w113, c0_n0_w114, c0_n0_w115, c0_n0_w116, c0_n0_w117, c0_n0_w118, c0_n0_w119, c0_n0_w120, c0_n0_w121, c0_n0_w122, c0_n0_w123, c0_n0_w124, c0_n0_w125, c0_n0_w126, c0_n0_w127, c0_n0_w128, c0_n0_w129, c0_n0_w130, c0_n0_w131, c0_n0_w132, c0_n0_w133, c0_n0_w134, c0_n0_w135, c0_n0_w136, c0_n0_w137, c0_n0_w138, c0_n0_w139, c0_n0_w140, c0_n0_w141, c0_n0_w142, c0_n0_w143, c0_n0_w144, c0_n0_w145, c0_n0_w146, c0_n0_w147, c0_n0_w148, c0_n0_w149, c0_n0_w150, c0_n0_w151, c0_n0_w152, c0_n0_w153, c0_n0_w154, c0_n0_w155, c0_n0_w156, c0_n0_w157, c0_n0_w158, c0_n0_w159, c0_n0_w160, c0_n0_w161, c0_n0_w162, c0_n0_w163, c0_n0_w164, c0_n0_w165, c0_n0_w166, c0_n0_w167, c0_n0_w168, c0_n0_w169, c0_n0_w170, c0_n0_w171, c0_n0_w172, c0_n0_w173, c0_n0_w174, c0_n0_w175, c0_n0_w176, c0_n0_w177, c0_n0_w178, c0_n0_w179, c0_n0_w180, c0_n0_w181, c0_n0_w182, c0_n0_w183, c0_n0_w184, c0_n0_w185, c0_n0_w186, c0_n0_w187, c0_n0_w188, c0_n0_w189, c0_n0_w190, c0_n0_w191, c0_n0_w192, c0_n0_w193, c0_n0_w194, c0_n0_w195, c0_n0_w196, c0_n0_w197, c0_n0_w198, c0_n0_w199, c0_n0_w200, c0_n1_w1, c0_n1_w2, c0_n1_w3, c0_n1_w4, c0_n1_w5, c0_n1_w6, c0_n1_w7, c0_n1_w8, c0_n1_w9, c0_n1_w10, c0_n1_w11, c0_n1_w12, c0_n1_w13, c0_n1_w14, c0_n1_w15, c0_n1_w16, c0_n1_w17, c0_n1_w18, c0_n1_w19, c0_n1_w20, c0_n1_w21, c0_n1_w22, c0_n1_w23, c0_n1_w24, c0_n1_w25, c0_n1_w26, c0_n1_w27, c0_n1_w28, c0_n1_w29, c0_n1_w30, c0_n1_w31, c0_n1_w32, c0_n1_w33, c0_n1_w34, c0_n1_w35, c0_n1_w36, c0_n1_w37, c0_n1_w38, c0_n1_w39, c0_n1_w40, c0_n1_w41, c0_n1_w42, c0_n1_w43, c0_n1_w44, c0_n1_w45, c0_n1_w46, c0_n1_w47, c0_n1_w48, c0_n1_w49, c0_n1_w50, c0_n1_w51, c0_n1_w52, c0_n1_w53, c0_n1_w54, c0_n1_w55, c0_n1_w56, c0_n1_w57, c0_n1_w58, c0_n1_w59, c0_n1_w60, c0_n1_w61, c0_n1_w62, c0_n1_w63, c0_n1_w64, c0_n1_w65, c0_n1_w66, c0_n1_w67, c0_n1_w68, c0_n1_w69, c0_n1_w70, c0_n1_w71, c0_n1_w72, c0_n1_w73, c0_n1_w74, c0_n1_w75, c0_n1_w76, c0_n1_w77, c0_n1_w78, c0_n1_w79, c0_n1_w80, c0_n1_w81, c0_n1_w82, c0_n1_w83, c0_n1_w84, c0_n1_w85, c0_n1_w86, c0_n1_w87, c0_n1_w88, c0_n1_w89, c0_n1_w90, c0_n1_w91, c0_n1_w92, c0_n1_w93, c0_n1_w94, c0_n1_w95, c0_n1_w96, c0_n1_w97, c0_n1_w98, c0_n1_w99, c0_n1_w100, c0_n1_w101, c0_n1_w102, c0_n1_w103, c0_n1_w104, c0_n1_w105, c0_n1_w106, c0_n1_w107, c0_n1_w108, c0_n1_w109, c0_n1_w110, c0_n1_w111, c0_n1_w112, c0_n1_w113, c0_n1_w114, c0_n1_w115, c0_n1_w116, c0_n1_w117, c0_n1_w118, c0_n1_w119, c0_n1_w120, c0_n1_w121, c0_n1_w122, c0_n1_w123, c0_n1_w124, c0_n1_w125, c0_n1_w126, c0_n1_w127, c0_n1_w128, c0_n1_w129, c0_n1_w130, c0_n1_w131, c0_n1_w132, c0_n1_w133, c0_n1_w134, c0_n1_w135, c0_n1_w136, c0_n1_w137, c0_n1_w138, c0_n1_w139, c0_n1_w140, c0_n1_w141, c0_n1_w142, c0_n1_w143, c0_n1_w144, c0_n1_w145, c0_n1_w146, c0_n1_w147, c0_n1_w148, c0_n1_w149, c0_n1_w150, c0_n1_w151, c0_n1_w152, c0_n1_w153, c0_n1_w154, c0_n1_w155, c0_n1_w156, c0_n1_w157, c0_n1_w158, c0_n1_w159, c0_n1_w160, c0_n1_w161, c0_n1_w162, c0_n1_w163, c0_n1_w164, c0_n1_w165, c0_n1_w166, c0_n1_w167, c0_n1_w168, c0_n1_w169, c0_n1_w170, c0_n1_w171, c0_n1_w172, c0_n1_w173, c0_n1_w174, c0_n1_w175, c0_n1_w176, c0_n1_w177, c0_n1_w178, c0_n1_w179, c0_n1_w180, c0_n1_w181, c0_n1_w182, c0_n1_w183, c0_n1_w184, c0_n1_w185, c0_n1_w186, c0_n1_w187, c0_n1_w188, c0_n1_w189, c0_n1_w190, c0_n1_w191, c0_n1_w192, c0_n1_w193, c0_n1_w194, c0_n1_w195, c0_n1_w196, c0_n1_w197, c0_n1_w198, c0_n1_w199, c0_n1_w200, c0_n2_w1, c0_n2_w2, c0_n2_w3, c0_n2_w4, c0_n2_w5, c0_n2_w6, c0_n2_w7, c0_n2_w8, c0_n2_w9, c0_n2_w10, c0_n2_w11, c0_n2_w12, c0_n2_w13, c0_n2_w14, c0_n2_w15, c0_n2_w16, c0_n2_w17, c0_n2_w18, c0_n2_w19, c0_n2_w20, c0_n2_w21, c0_n2_w22, c0_n2_w23, c0_n2_w24, c0_n2_w25, c0_n2_w26, c0_n2_w27, c0_n2_w28, c0_n2_w29, c0_n2_w30, c0_n2_w31, c0_n2_w32, c0_n2_w33, c0_n2_w34, c0_n2_w35, c0_n2_w36, c0_n2_w37, c0_n2_w38, c0_n2_w39, c0_n2_w40, c0_n2_w41, c0_n2_w42, c0_n2_w43, c0_n2_w44, c0_n2_w45, c0_n2_w46, c0_n2_w47, c0_n2_w48, c0_n2_w49, c0_n2_w50, c0_n2_w51, c0_n2_w52, c0_n2_w53, c0_n2_w54, c0_n2_w55, c0_n2_w56, c0_n2_w57, c0_n2_w58, c0_n2_w59, c0_n2_w60, c0_n2_w61, c0_n2_w62, c0_n2_w63, c0_n2_w64, c0_n2_w65, c0_n2_w66, c0_n2_w67, c0_n2_w68, c0_n2_w69, c0_n2_w70, c0_n2_w71, c0_n2_w72, c0_n2_w73, c0_n2_w74, c0_n2_w75, c0_n2_w76, c0_n2_w77, c0_n2_w78, c0_n2_w79, c0_n2_w80, c0_n2_w81, c0_n2_w82, c0_n2_w83, c0_n2_w84, c0_n2_w85, c0_n2_w86, c0_n2_w87, c0_n2_w88, c0_n2_w89, c0_n2_w90, c0_n2_w91, c0_n2_w92, c0_n2_w93, c0_n2_w94, c0_n2_w95, c0_n2_w96, c0_n2_w97, c0_n2_w98, c0_n2_w99, c0_n2_w100, c0_n2_w101, c0_n2_w102, c0_n2_w103, c0_n2_w104, c0_n2_w105, c0_n2_w106, c0_n2_w107, c0_n2_w108, c0_n2_w109, c0_n2_w110, c0_n2_w111, c0_n2_w112, c0_n2_w113, c0_n2_w114, c0_n2_w115, c0_n2_w116, c0_n2_w117, c0_n2_w118, c0_n2_w119, c0_n2_w120, c0_n2_w121, c0_n2_w122, c0_n2_w123, c0_n2_w124, c0_n2_w125, c0_n2_w126, c0_n2_w127, c0_n2_w128, c0_n2_w129, c0_n2_w130, c0_n2_w131, c0_n2_w132, c0_n2_w133, c0_n2_w134, c0_n2_w135, c0_n2_w136, c0_n2_w137, c0_n2_w138, c0_n2_w139, c0_n2_w140, c0_n2_w141, c0_n2_w142, c0_n2_w143, c0_n2_w144, c0_n2_w145, c0_n2_w146, c0_n2_w147, c0_n2_w148, c0_n2_w149, c0_n2_w150, c0_n2_w151, c0_n2_w152, c0_n2_w153, c0_n2_w154, c0_n2_w155, c0_n2_w156, c0_n2_w157, c0_n2_w158, c0_n2_w159, c0_n2_w160, c0_n2_w161, c0_n2_w162, c0_n2_w163, c0_n2_w164, c0_n2_w165, c0_n2_w166, c0_n2_w167, c0_n2_w168, c0_n2_w169, c0_n2_w170, c0_n2_w171, c0_n2_w172, c0_n2_w173, c0_n2_w174, c0_n2_w175, c0_n2_w176, c0_n2_w177, c0_n2_w178, c0_n2_w179, c0_n2_w180, c0_n2_w181, c0_n2_w182, c0_n2_w183, c0_n2_w184, c0_n2_w185, c0_n2_w186, c0_n2_w187, c0_n2_w188, c0_n2_w189, c0_n2_w190, c0_n2_w191, c0_n2_w192, c0_n2_w193, c0_n2_w194, c0_n2_w195, c0_n2_w196, c0_n2_w197, c0_n2_w198, c0_n2_w199, c0_n2_w200, c0_n3_w1, c0_n3_w2, c0_n3_w3, c0_n3_w4, c0_n3_w5, c0_n3_w6, c0_n3_w7, c0_n3_w8, c0_n3_w9, c0_n3_w10, c0_n3_w11, c0_n3_w12, c0_n3_w13, c0_n3_w14, c0_n3_w15, c0_n3_w16, c0_n3_w17, c0_n3_w18, c0_n3_w19, c0_n3_w20, c0_n3_w21, c0_n3_w22, c0_n3_w23, c0_n3_w24, c0_n3_w25, c0_n3_w26, c0_n3_w27, c0_n3_w28, c0_n3_w29, c0_n3_w30, c0_n3_w31, c0_n3_w32, c0_n3_w33, c0_n3_w34, c0_n3_w35, c0_n3_w36, c0_n3_w37, c0_n3_w38, c0_n3_w39, c0_n3_w40, c0_n3_w41, c0_n3_w42, c0_n3_w43, c0_n3_w44, c0_n3_w45, c0_n3_w46, c0_n3_w47, c0_n3_w48, c0_n3_w49, c0_n3_w50, c0_n3_w51, c0_n3_w52, c0_n3_w53, c0_n3_w54, c0_n3_w55, c0_n3_w56, c0_n3_w57, c0_n3_w58, c0_n3_w59, c0_n3_w60, c0_n3_w61, c0_n3_w62, c0_n3_w63, c0_n3_w64, c0_n3_w65, c0_n3_w66, c0_n3_w67, c0_n3_w68, c0_n3_w69, c0_n3_w70, c0_n3_w71, c0_n3_w72, c0_n3_w73, c0_n3_w74, c0_n3_w75, c0_n3_w76, c0_n3_w77, c0_n3_w78, c0_n3_w79, c0_n3_w80, c0_n3_w81, c0_n3_w82, c0_n3_w83, c0_n3_w84, c0_n3_w85, c0_n3_w86, c0_n3_w87, c0_n3_w88, c0_n3_w89, c0_n3_w90, c0_n3_w91, c0_n3_w92, c0_n3_w93, c0_n3_w94, c0_n3_w95, c0_n3_w96, c0_n3_w97, c0_n3_w98, c0_n3_w99, c0_n3_w100, c0_n3_w101, c0_n3_w102, c0_n3_w103, c0_n3_w104, c0_n3_w105, c0_n3_w106, c0_n3_w107, c0_n3_w108, c0_n3_w109, c0_n3_w110, c0_n3_w111, c0_n3_w112, c0_n3_w113, c0_n3_w114, c0_n3_w115, c0_n3_w116, c0_n3_w117, c0_n3_w118, c0_n3_w119, c0_n3_w120, c0_n3_w121, c0_n3_w122, c0_n3_w123, c0_n3_w124, c0_n3_w125, c0_n3_w126, c0_n3_w127, c0_n3_w128, c0_n3_w129, c0_n3_w130, c0_n3_w131, c0_n3_w132, c0_n3_w133, c0_n3_w134, c0_n3_w135, c0_n3_w136, c0_n3_w137, c0_n3_w138, c0_n3_w139, c0_n3_w140, c0_n3_w141, c0_n3_w142, c0_n3_w143, c0_n3_w144, c0_n3_w145, c0_n3_w146, c0_n3_w147, c0_n3_w148, c0_n3_w149, c0_n3_w150, c0_n3_w151, c0_n3_w152, c0_n3_w153, c0_n3_w154, c0_n3_w155, c0_n3_w156, c0_n3_w157, c0_n3_w158, c0_n3_w159, c0_n3_w160, c0_n3_w161, c0_n3_w162, c0_n3_w163, c0_n3_w164, c0_n3_w165, c0_n3_w166, c0_n3_w167, c0_n3_w168, c0_n3_w169, c0_n3_w170, c0_n3_w171, c0_n3_w172, c0_n3_w173, c0_n3_w174, c0_n3_w175, c0_n3_w176, c0_n3_w177, c0_n3_w178, c0_n3_w179, c0_n3_w180, c0_n3_w181, c0_n3_w182, c0_n3_w183, c0_n3_w184, c0_n3_w185, c0_n3_w186, c0_n3_w187, c0_n3_w188, c0_n3_w189, c0_n3_w190, c0_n3_w191, c0_n3_w192, c0_n3_w193, c0_n3_w194, c0_n3_w195, c0_n3_w196, c0_n3_w197, c0_n3_w198, c0_n3_w199, c0_n3_w200, c0_n4_w1, c0_n4_w2, c0_n4_w3, c0_n4_w4, c0_n4_w5, c0_n4_w6, c0_n4_w7, c0_n4_w8, c0_n4_w9, c0_n4_w10, c0_n4_w11, c0_n4_w12, c0_n4_w13, c0_n4_w14, c0_n4_w15, c0_n4_w16, c0_n4_w17, c0_n4_w18, c0_n4_w19, c0_n4_w20, c0_n4_w21, c0_n4_w22, c0_n4_w23, c0_n4_w24, c0_n4_w25, c0_n4_w26, c0_n4_w27, c0_n4_w28, c0_n4_w29, c0_n4_w30, c0_n4_w31, c0_n4_w32, c0_n4_w33, c0_n4_w34, c0_n4_w35, c0_n4_w36, c0_n4_w37, c0_n4_w38, c0_n4_w39, c0_n4_w40, c0_n4_w41, c0_n4_w42, c0_n4_w43, c0_n4_w44, c0_n4_w45, c0_n4_w46, c0_n4_w47, c0_n4_w48, c0_n4_w49, c0_n4_w50, c0_n4_w51, c0_n4_w52, c0_n4_w53, c0_n4_w54, c0_n4_w55, c0_n4_w56, c0_n4_w57, c0_n4_w58, c0_n4_w59, c0_n4_w60, c0_n4_w61, c0_n4_w62, c0_n4_w63, c0_n4_w64, c0_n4_w65, c0_n4_w66, c0_n4_w67, c0_n4_w68, c0_n4_w69, c0_n4_w70, c0_n4_w71, c0_n4_w72, c0_n4_w73, c0_n4_w74, c0_n4_w75, c0_n4_w76, c0_n4_w77, c0_n4_w78, c0_n4_w79, c0_n4_w80, c0_n4_w81, c0_n4_w82, c0_n4_w83, c0_n4_w84, c0_n4_w85, c0_n4_w86, c0_n4_w87, c0_n4_w88, c0_n4_w89, c0_n4_w90, c0_n4_w91, c0_n4_w92, c0_n4_w93, c0_n4_w94, c0_n4_w95, c0_n4_w96, c0_n4_w97, c0_n4_w98, c0_n4_w99, c0_n4_w100, c0_n4_w101, c0_n4_w102, c0_n4_w103, c0_n4_w104, c0_n4_w105, c0_n4_w106, c0_n4_w107, c0_n4_w108, c0_n4_w109, c0_n4_w110, c0_n4_w111, c0_n4_w112, c0_n4_w113, c0_n4_w114, c0_n4_w115, c0_n4_w116, c0_n4_w117, c0_n4_w118, c0_n4_w119, c0_n4_w120, c0_n4_w121, c0_n4_w122, c0_n4_w123, c0_n4_w124, c0_n4_w125, c0_n4_w126, c0_n4_w127, c0_n4_w128, c0_n4_w129, c0_n4_w130, c0_n4_w131, c0_n4_w132, c0_n4_w133, c0_n4_w134, c0_n4_w135, c0_n4_w136, c0_n4_w137, c0_n4_w138, c0_n4_w139, c0_n4_w140, c0_n4_w141, c0_n4_w142, c0_n4_w143, c0_n4_w144, c0_n4_w145, c0_n4_w146, c0_n4_w147, c0_n4_w148, c0_n4_w149, c0_n4_w150, c0_n4_w151, c0_n4_w152, c0_n4_w153, c0_n4_w154, c0_n4_w155, c0_n4_w156, c0_n4_w157, c0_n4_w158, c0_n4_w159, c0_n4_w160, c0_n4_w161, c0_n4_w162, c0_n4_w163, c0_n4_w164, c0_n4_w165, c0_n4_w166, c0_n4_w167, c0_n4_w168, c0_n4_w169, c0_n4_w170, c0_n4_w171, c0_n4_w172, c0_n4_w173, c0_n4_w174, c0_n4_w175, c0_n4_w176, c0_n4_w177, c0_n4_w178, c0_n4_w179, c0_n4_w180, c0_n4_w181, c0_n4_w182, c0_n4_w183, c0_n4_w184, c0_n4_w185, c0_n4_w186, c0_n4_w187, c0_n4_w188, c0_n4_w189, c0_n4_w190, c0_n4_w191, c0_n4_w192, c0_n4_w193, c0_n4_w194, c0_n4_w195, c0_n4_w196, c0_n4_w197, c0_n4_w198, c0_n4_w199, c0_n4_w200, c0_n5_w1, c0_n5_w2, c0_n5_w3, c0_n5_w4, c0_n5_w5, c0_n5_w6, c0_n5_w7, c0_n5_w8, c0_n5_w9, c0_n5_w10, c0_n5_w11, c0_n5_w12, c0_n5_w13, c0_n5_w14, c0_n5_w15, c0_n5_w16, c0_n5_w17, c0_n5_w18, c0_n5_w19, c0_n5_w20, c0_n5_w21, c0_n5_w22, c0_n5_w23, c0_n5_w24, c0_n5_w25, c0_n5_w26, c0_n5_w27, c0_n5_w28, c0_n5_w29, c0_n5_w30, c0_n5_w31, c0_n5_w32, c0_n5_w33, c0_n5_w34, c0_n5_w35, c0_n5_w36, c0_n5_w37, c0_n5_w38, c0_n5_w39, c0_n5_w40, c0_n5_w41, c0_n5_w42, c0_n5_w43, c0_n5_w44, c0_n5_w45, c0_n5_w46, c0_n5_w47, c0_n5_w48, c0_n5_w49, c0_n5_w50, c0_n5_w51, c0_n5_w52, c0_n5_w53, c0_n5_w54, c0_n5_w55, c0_n5_w56, c0_n5_w57, c0_n5_w58, c0_n5_w59, c0_n5_w60, c0_n5_w61, c0_n5_w62, c0_n5_w63, c0_n5_w64, c0_n5_w65, c0_n5_w66, c0_n5_w67, c0_n5_w68, c0_n5_w69, c0_n5_w70, c0_n5_w71, c0_n5_w72, c0_n5_w73, c0_n5_w74, c0_n5_w75, c0_n5_w76, c0_n5_w77, c0_n5_w78, c0_n5_w79, c0_n5_w80, c0_n5_w81, c0_n5_w82, c0_n5_w83, c0_n5_w84, c0_n5_w85, c0_n5_w86, c0_n5_w87, c0_n5_w88, c0_n5_w89, c0_n5_w90, c0_n5_w91, c0_n5_w92, c0_n5_w93, c0_n5_w94, c0_n5_w95, c0_n5_w96, c0_n5_w97, c0_n5_w98, c0_n5_w99, c0_n5_w100, c0_n5_w101, c0_n5_w102, c0_n5_w103, c0_n5_w104, c0_n5_w105, c0_n5_w106, c0_n5_w107, c0_n5_w108, c0_n5_w109, c0_n5_w110, c0_n5_w111, c0_n5_w112, c0_n5_w113, c0_n5_w114, c0_n5_w115, c0_n5_w116, c0_n5_w117, c0_n5_w118, c0_n5_w119, c0_n5_w120, c0_n5_w121, c0_n5_w122, c0_n5_w123, c0_n5_w124, c0_n5_w125, c0_n5_w126, c0_n5_w127, c0_n5_w128, c0_n5_w129, c0_n5_w130, c0_n5_w131, c0_n5_w132, c0_n5_w133, c0_n5_w134, c0_n5_w135, c0_n5_w136, c0_n5_w137, c0_n5_w138, c0_n5_w139, c0_n5_w140, c0_n5_w141, c0_n5_w142, c0_n5_w143, c0_n5_w144, c0_n5_w145, c0_n5_w146, c0_n5_w147, c0_n5_w148, c0_n5_w149, c0_n5_w150, c0_n5_w151, c0_n5_w152, c0_n5_w153, c0_n5_w154, c0_n5_w155, c0_n5_w156, c0_n5_w157, c0_n5_w158, c0_n5_w159, c0_n5_w160, c0_n5_w161, c0_n5_w162, c0_n5_w163, c0_n5_w164, c0_n5_w165, c0_n5_w166, c0_n5_w167, c0_n5_w168, c0_n5_w169, c0_n5_w170, c0_n5_w171, c0_n5_w172, c0_n5_w173, c0_n5_w174, c0_n5_w175, c0_n5_w176, c0_n5_w177, c0_n5_w178, c0_n5_w179, c0_n5_w180, c0_n5_w181, c0_n5_w182, c0_n5_w183, c0_n5_w184, c0_n5_w185, c0_n5_w186, c0_n5_w187, c0_n5_w188, c0_n5_w189, c0_n5_w190, c0_n5_w191, c0_n5_w192, c0_n5_w193, c0_n5_w194, c0_n5_w195, c0_n5_w196, c0_n5_w197, c0_n5_w198, c0_n5_w199, c0_n5_w200, c0_n6_w1, c0_n6_w2, c0_n6_w3, c0_n6_w4, c0_n6_w5, c0_n6_w6, c0_n6_w7, c0_n6_w8, c0_n6_w9, c0_n6_w10, c0_n6_w11, c0_n6_w12, c0_n6_w13, c0_n6_w14, c0_n6_w15, c0_n6_w16, c0_n6_w17, c0_n6_w18, c0_n6_w19, c0_n6_w20, c0_n6_w21, c0_n6_w22, c0_n6_w23, c0_n6_w24, c0_n6_w25, c0_n6_w26, c0_n6_w27, c0_n6_w28, c0_n6_w29, c0_n6_w30, c0_n6_w31, c0_n6_w32, c0_n6_w33, c0_n6_w34, c0_n6_w35, c0_n6_w36, c0_n6_w37, c0_n6_w38, c0_n6_w39, c0_n6_w40, c0_n6_w41, c0_n6_w42, c0_n6_w43, c0_n6_w44, c0_n6_w45, c0_n6_w46, c0_n6_w47, c0_n6_w48, c0_n6_w49, c0_n6_w50, c0_n6_w51, c0_n6_w52, c0_n6_w53, c0_n6_w54, c0_n6_w55, c0_n6_w56, c0_n6_w57, c0_n6_w58, c0_n6_w59, c0_n6_w60, c0_n6_w61, c0_n6_w62, c0_n6_w63, c0_n6_w64, c0_n6_w65, c0_n6_w66, c0_n6_w67, c0_n6_w68, c0_n6_w69, c0_n6_w70, c0_n6_w71, c0_n6_w72, c0_n6_w73, c0_n6_w74, c0_n6_w75, c0_n6_w76, c0_n6_w77, c0_n6_w78, c0_n6_w79, c0_n6_w80, c0_n6_w81, c0_n6_w82, c0_n6_w83, c0_n6_w84, c0_n6_w85, c0_n6_w86, c0_n6_w87, c0_n6_w88, c0_n6_w89, c0_n6_w90, c0_n6_w91, c0_n6_w92, c0_n6_w93, c0_n6_w94, c0_n6_w95, c0_n6_w96, c0_n6_w97, c0_n6_w98, c0_n6_w99, c0_n6_w100, c0_n6_w101, c0_n6_w102, c0_n6_w103, c0_n6_w104, c0_n6_w105, c0_n6_w106, c0_n6_w107, c0_n6_w108, c0_n6_w109, c0_n6_w110, c0_n6_w111, c0_n6_w112, c0_n6_w113, c0_n6_w114, c0_n6_w115, c0_n6_w116, c0_n6_w117, c0_n6_w118, c0_n6_w119, c0_n6_w120, c0_n6_w121, c0_n6_w122, c0_n6_w123, c0_n6_w124, c0_n6_w125, c0_n6_w126, c0_n6_w127, c0_n6_w128, c0_n6_w129, c0_n6_w130, c0_n6_w131, c0_n6_w132, c0_n6_w133, c0_n6_w134, c0_n6_w135, c0_n6_w136, c0_n6_w137, c0_n6_w138, c0_n6_w139, c0_n6_w140, c0_n6_w141, c0_n6_w142, c0_n6_w143, c0_n6_w144, c0_n6_w145, c0_n6_w146, c0_n6_w147, c0_n6_w148, c0_n6_w149, c0_n6_w150, c0_n6_w151, c0_n6_w152, c0_n6_w153, c0_n6_w154, c0_n6_w155, c0_n6_w156, c0_n6_w157, c0_n6_w158, c0_n6_w159, c0_n6_w160, c0_n6_w161, c0_n6_w162, c0_n6_w163, c0_n6_w164, c0_n6_w165, c0_n6_w166, c0_n6_w167, c0_n6_w168, c0_n6_w169, c0_n6_w170, c0_n6_w171, c0_n6_w172, c0_n6_w173, c0_n6_w174, c0_n6_w175, c0_n6_w176, c0_n6_w177, c0_n6_w178, c0_n6_w179, c0_n6_w180, c0_n6_w181, c0_n6_w182, c0_n6_w183, c0_n6_w184, c0_n6_w185, c0_n6_w186, c0_n6_w187, c0_n6_w188, c0_n6_w189, c0_n6_w190, c0_n6_w191, c0_n6_w192, c0_n6_w193, c0_n6_w194, c0_n6_w195, c0_n6_w196, c0_n6_w197, c0_n6_w198, c0_n6_w199, c0_n6_w200, c0_n7_w1, c0_n7_w2, c0_n7_w3, c0_n7_w4, c0_n7_w5, c0_n7_w6, c0_n7_w7, c0_n7_w8, c0_n7_w9, c0_n7_w10, c0_n7_w11, c0_n7_w12, c0_n7_w13, c0_n7_w14, c0_n7_w15, c0_n7_w16, c0_n7_w17, c0_n7_w18, c0_n7_w19, c0_n7_w20, c0_n7_w21, c0_n7_w22, c0_n7_w23, c0_n7_w24, c0_n7_w25, c0_n7_w26, c0_n7_w27, c0_n7_w28, c0_n7_w29, c0_n7_w30, c0_n7_w31, c0_n7_w32, c0_n7_w33, c0_n7_w34, c0_n7_w35, c0_n7_w36, c0_n7_w37, c0_n7_w38, c0_n7_w39, c0_n7_w40, c0_n7_w41, c0_n7_w42, c0_n7_w43, c0_n7_w44, c0_n7_w45, c0_n7_w46, c0_n7_w47, c0_n7_w48, c0_n7_w49, c0_n7_w50, c0_n7_w51, c0_n7_w52, c0_n7_w53, c0_n7_w54, c0_n7_w55, c0_n7_w56, c0_n7_w57, c0_n7_w58, c0_n7_w59, c0_n7_w60, c0_n7_w61, c0_n7_w62, c0_n7_w63, c0_n7_w64, c0_n7_w65, c0_n7_w66, c0_n7_w67, c0_n7_w68, c0_n7_w69, c0_n7_w70, c0_n7_w71, c0_n7_w72, c0_n7_w73, c0_n7_w74, c0_n7_w75, c0_n7_w76, c0_n7_w77, c0_n7_w78, c0_n7_w79, c0_n7_w80, c0_n7_w81, c0_n7_w82, c0_n7_w83, c0_n7_w84, c0_n7_w85, c0_n7_w86, c0_n7_w87, c0_n7_w88, c0_n7_w89, c0_n7_w90, c0_n7_w91, c0_n7_w92, c0_n7_w93, c0_n7_w94, c0_n7_w95, c0_n7_w96, c0_n7_w97, c0_n7_w98, c0_n7_w99, c0_n7_w100, c0_n7_w101, c0_n7_w102, c0_n7_w103, c0_n7_w104, c0_n7_w105, c0_n7_w106, c0_n7_w107, c0_n7_w108, c0_n7_w109, c0_n7_w110, c0_n7_w111, c0_n7_w112, c0_n7_w113, c0_n7_w114, c0_n7_w115, c0_n7_w116, c0_n7_w117, c0_n7_w118, c0_n7_w119, c0_n7_w120, c0_n7_w121, c0_n7_w122, c0_n7_w123, c0_n7_w124, c0_n7_w125, c0_n7_w126, c0_n7_w127, c0_n7_w128, c0_n7_w129, c0_n7_w130, c0_n7_w131, c0_n7_w132, c0_n7_w133, c0_n7_w134, c0_n7_w135, c0_n7_w136, c0_n7_w137, c0_n7_w138, c0_n7_w139, c0_n7_w140, c0_n7_w141, c0_n7_w142, c0_n7_w143, c0_n7_w144, c0_n7_w145, c0_n7_w146, c0_n7_w147, c0_n7_w148, c0_n7_w149, c0_n7_w150, c0_n7_w151, c0_n7_w152, c0_n7_w153, c0_n7_w154, c0_n7_w155, c0_n7_w156, c0_n7_w157, c0_n7_w158, c0_n7_w159, c0_n7_w160, c0_n7_w161, c0_n7_w162, c0_n7_w163, c0_n7_w164, c0_n7_w165, c0_n7_w166, c0_n7_w167, c0_n7_w168, c0_n7_w169, c0_n7_w170, c0_n7_w171, c0_n7_w172, c0_n7_w173, c0_n7_w174, c0_n7_w175, c0_n7_w176, c0_n7_w177, c0_n7_w178, c0_n7_w179, c0_n7_w180, c0_n7_w181, c0_n7_w182, c0_n7_w183, c0_n7_w184, c0_n7_w185, c0_n7_w186, c0_n7_w187, c0_n7_w188, c0_n7_w189, c0_n7_w190, c0_n7_w191, c0_n7_w192, c0_n7_w193, c0_n7_w194, c0_n7_w195, c0_n7_w196, c0_n7_w197, c0_n7_w198, c0_n7_w199, c0_n7_w200, c0_n8_w1, c0_n8_w2, c0_n8_w3, c0_n8_w4, c0_n8_w5, c0_n8_w6, c0_n8_w7, c0_n8_w8, c0_n8_w9, c0_n8_w10, c0_n8_w11, c0_n8_w12, c0_n8_w13, c0_n8_w14, c0_n8_w15, c0_n8_w16, c0_n8_w17, c0_n8_w18, c0_n8_w19, c0_n8_w20, c0_n8_w21, c0_n8_w22, c0_n8_w23, c0_n8_w24, c0_n8_w25, c0_n8_w26, c0_n8_w27, c0_n8_w28, c0_n8_w29, c0_n8_w30, c0_n8_w31, c0_n8_w32, c0_n8_w33, c0_n8_w34, c0_n8_w35, c0_n8_w36, c0_n8_w37, c0_n8_w38, c0_n8_w39, c0_n8_w40, c0_n8_w41, c0_n8_w42, c0_n8_w43, c0_n8_w44, c0_n8_w45, c0_n8_w46, c0_n8_w47, c0_n8_w48, c0_n8_w49, c0_n8_w50, c0_n8_w51, c0_n8_w52, c0_n8_w53, c0_n8_w54, c0_n8_w55, c0_n8_w56, c0_n8_w57, c0_n8_w58, c0_n8_w59, c0_n8_w60, c0_n8_w61, c0_n8_w62, c0_n8_w63, c0_n8_w64, c0_n8_w65, c0_n8_w66, c0_n8_w67, c0_n8_w68, c0_n8_w69, c0_n8_w70, c0_n8_w71, c0_n8_w72, c0_n8_w73, c0_n8_w74, c0_n8_w75, c0_n8_w76, c0_n8_w77, c0_n8_w78, c0_n8_w79, c0_n8_w80, c0_n8_w81, c0_n8_w82, c0_n8_w83, c0_n8_w84, c0_n8_w85, c0_n8_w86, c0_n8_w87, c0_n8_w88, c0_n8_w89, c0_n8_w90, c0_n8_w91, c0_n8_w92, c0_n8_w93, c0_n8_w94, c0_n8_w95, c0_n8_w96, c0_n8_w97, c0_n8_w98, c0_n8_w99, c0_n8_w100, c0_n8_w101, c0_n8_w102, c0_n8_w103, c0_n8_w104, c0_n8_w105, c0_n8_w106, c0_n8_w107, c0_n8_w108, c0_n8_w109, c0_n8_w110, c0_n8_w111, c0_n8_w112, c0_n8_w113, c0_n8_w114, c0_n8_w115, c0_n8_w116, c0_n8_w117, c0_n8_w118, c0_n8_w119, c0_n8_w120, c0_n8_w121, c0_n8_w122, c0_n8_w123, c0_n8_w124, c0_n8_w125, c0_n8_w126, c0_n8_w127, c0_n8_w128, c0_n8_w129, c0_n8_w130, c0_n8_w131, c0_n8_w132, c0_n8_w133, c0_n8_w134, c0_n8_w135, c0_n8_w136, c0_n8_w137, c0_n8_w138, c0_n8_w139, c0_n8_w140, c0_n8_w141, c0_n8_w142, c0_n8_w143, c0_n8_w144, c0_n8_w145, c0_n8_w146, c0_n8_w147, c0_n8_w148, c0_n8_w149, c0_n8_w150, c0_n8_w151, c0_n8_w152, c0_n8_w153, c0_n8_w154, c0_n8_w155, c0_n8_w156, c0_n8_w157, c0_n8_w158, c0_n8_w159, c0_n8_w160, c0_n8_w161, c0_n8_w162, c0_n8_w163, c0_n8_w164, c0_n8_w165, c0_n8_w166, c0_n8_w167, c0_n8_w168, c0_n8_w169, c0_n8_w170, c0_n8_w171, c0_n8_w172, c0_n8_w173, c0_n8_w174, c0_n8_w175, c0_n8_w176, c0_n8_w177, c0_n8_w178, c0_n8_w179, c0_n8_w180, c0_n8_w181, c0_n8_w182, c0_n8_w183, c0_n8_w184, c0_n8_w185, c0_n8_w186, c0_n8_w187, c0_n8_w188, c0_n8_w189, c0_n8_w190, c0_n8_w191, c0_n8_w192, c0_n8_w193, c0_n8_w194, c0_n8_w195, c0_n8_w196, c0_n8_w197, c0_n8_w198, c0_n8_w199, c0_n8_w200, c0_n9_w1, c0_n9_w2, c0_n9_w3, c0_n9_w4, c0_n9_w5, c0_n9_w6, c0_n9_w7, c0_n9_w8, c0_n9_w9, c0_n9_w10, c0_n9_w11, c0_n9_w12, c0_n9_w13, c0_n9_w14, c0_n9_w15, c0_n9_w16, c0_n9_w17, c0_n9_w18, c0_n9_w19, c0_n9_w20, c0_n9_w21, c0_n9_w22, c0_n9_w23, c0_n9_w24, c0_n9_w25, c0_n9_w26, c0_n9_w27, c0_n9_w28, c0_n9_w29, c0_n9_w30, c0_n9_w31, c0_n9_w32, c0_n9_w33, c0_n9_w34, c0_n9_w35, c0_n9_w36, c0_n9_w37, c0_n9_w38, c0_n9_w39, c0_n9_w40, c0_n9_w41, c0_n9_w42, c0_n9_w43, c0_n9_w44, c0_n9_w45, c0_n9_w46, c0_n9_w47, c0_n9_w48, c0_n9_w49, c0_n9_w50, c0_n9_w51, c0_n9_w52, c0_n9_w53, c0_n9_w54, c0_n9_w55, c0_n9_w56, c0_n9_w57, c0_n9_w58, c0_n9_w59, c0_n9_w60, c0_n9_w61, c0_n9_w62, c0_n9_w63, c0_n9_w64, c0_n9_w65, c0_n9_w66, c0_n9_w67, c0_n9_w68, c0_n9_w69, c0_n9_w70, c0_n9_w71, c0_n9_w72, c0_n9_w73, c0_n9_w74, c0_n9_w75, c0_n9_w76, c0_n9_w77, c0_n9_w78, c0_n9_w79, c0_n9_w80, c0_n9_w81, c0_n9_w82, c0_n9_w83, c0_n9_w84, c0_n9_w85, c0_n9_w86, c0_n9_w87, c0_n9_w88, c0_n9_w89, c0_n9_w90, c0_n9_w91, c0_n9_w92, c0_n9_w93, c0_n9_w94, c0_n9_w95, c0_n9_w96, c0_n9_w97, c0_n9_w98, c0_n9_w99, c0_n9_w100, c0_n9_w101, c0_n9_w102, c0_n9_w103, c0_n9_w104, c0_n9_w105, c0_n9_w106, c0_n9_w107, c0_n9_w108, c0_n9_w109, c0_n9_w110, c0_n9_w111, c0_n9_w112, c0_n9_w113, c0_n9_w114, c0_n9_w115, c0_n9_w116, c0_n9_w117, c0_n9_w118, c0_n9_w119, c0_n9_w120, c0_n9_w121, c0_n9_w122, c0_n9_w123, c0_n9_w124, c0_n9_w125, c0_n9_w126, c0_n9_w127, c0_n9_w128, c0_n9_w129, c0_n9_w130, c0_n9_w131, c0_n9_w132, c0_n9_w133, c0_n9_w134, c0_n9_w135, c0_n9_w136, c0_n9_w137, c0_n9_w138, c0_n9_w139, c0_n9_w140, c0_n9_w141, c0_n9_w142, c0_n9_w143, c0_n9_w144, c0_n9_w145, c0_n9_w146, c0_n9_w147, c0_n9_w148, c0_n9_w149, c0_n9_w150, c0_n9_w151, c0_n9_w152, c0_n9_w153, c0_n9_w154, c0_n9_w155, c0_n9_w156, c0_n9_w157, c0_n9_w158, c0_n9_w159, c0_n9_w160, c0_n9_w161, c0_n9_w162, c0_n9_w163, c0_n9_w164, c0_n9_w165, c0_n9_w166, c0_n9_w167, c0_n9_w168, c0_n9_w169, c0_n9_w170, c0_n9_w171, c0_n9_w172, c0_n9_w173, c0_n9_w174, c0_n9_w175, c0_n9_w176, c0_n9_w177, c0_n9_w178, c0_n9_w179, c0_n9_w180, c0_n9_w181, c0_n9_w182, c0_n9_w183, c0_n9_w184, c0_n9_w185, c0_n9_w186, c0_n9_w187, c0_n9_w188, c0_n9_w189, c0_n9_w190, c0_n9_w191, c0_n9_w192, c0_n9_w193, c0_n9_w194, c0_n9_w195, c0_n9_w196, c0_n9_w197, c0_n9_w198, c0_n9_w199, c0_n9_w200, c0_n10_w1, c0_n10_w2, c0_n10_w3, c0_n10_w4, c0_n10_w5, c0_n10_w6, c0_n10_w7, c0_n10_w8, c0_n10_w9, c0_n10_w10, c0_n10_w11, c0_n10_w12, c0_n10_w13, c0_n10_w14, c0_n10_w15, c0_n10_w16, c0_n10_w17, c0_n10_w18, c0_n10_w19, c0_n10_w20, c0_n10_w21, c0_n10_w22, c0_n10_w23, c0_n10_w24, c0_n10_w25, c0_n10_w26, c0_n10_w27, c0_n10_w28, c0_n10_w29, c0_n10_w30, c0_n10_w31, c0_n10_w32, c0_n10_w33, c0_n10_w34, c0_n10_w35, c0_n10_w36, c0_n10_w37, c0_n10_w38, c0_n10_w39, c0_n10_w40, c0_n10_w41, c0_n10_w42, c0_n10_w43, c0_n10_w44, c0_n10_w45, c0_n10_w46, c0_n10_w47, c0_n10_w48, c0_n10_w49, c0_n10_w50, c0_n10_w51, c0_n10_w52, c0_n10_w53, c0_n10_w54, c0_n10_w55, c0_n10_w56, c0_n10_w57, c0_n10_w58, c0_n10_w59, c0_n10_w60, c0_n10_w61, c0_n10_w62, c0_n10_w63, c0_n10_w64, c0_n10_w65, c0_n10_w66, c0_n10_w67, c0_n10_w68, c0_n10_w69, c0_n10_w70, c0_n10_w71, c0_n10_w72, c0_n10_w73, c0_n10_w74, c0_n10_w75, c0_n10_w76, c0_n10_w77, c0_n10_w78, c0_n10_w79, c0_n10_w80, c0_n10_w81, c0_n10_w82, c0_n10_w83, c0_n10_w84, c0_n10_w85, c0_n10_w86, c0_n10_w87, c0_n10_w88, c0_n10_w89, c0_n10_w90, c0_n10_w91, c0_n10_w92, c0_n10_w93, c0_n10_w94, c0_n10_w95, c0_n10_w96, c0_n10_w97, c0_n10_w98, c0_n10_w99, c0_n10_w100, c0_n10_w101, c0_n10_w102, c0_n10_w103, c0_n10_w104, c0_n10_w105, c0_n10_w106, c0_n10_w107, c0_n10_w108, c0_n10_w109, c0_n10_w110, c0_n10_w111, c0_n10_w112, c0_n10_w113, c0_n10_w114, c0_n10_w115, c0_n10_w116, c0_n10_w117, c0_n10_w118, c0_n10_w119, c0_n10_w120, c0_n10_w121, c0_n10_w122, c0_n10_w123, c0_n10_w124, c0_n10_w125, c0_n10_w126, c0_n10_w127, c0_n10_w128, c0_n10_w129, c0_n10_w130, c0_n10_w131, c0_n10_w132, c0_n10_w133, c0_n10_w134, c0_n10_w135, c0_n10_w136, c0_n10_w137, c0_n10_w138, c0_n10_w139, c0_n10_w140, c0_n10_w141, c0_n10_w142, c0_n10_w143, c0_n10_w144, c0_n10_w145, c0_n10_w146, c0_n10_w147, c0_n10_w148, c0_n10_w149, c0_n10_w150, c0_n10_w151, c0_n10_w152, c0_n10_w153, c0_n10_w154, c0_n10_w155, c0_n10_w156, c0_n10_w157, c0_n10_w158, c0_n10_w159, c0_n10_w160, c0_n10_w161, c0_n10_w162, c0_n10_w163, c0_n10_w164, c0_n10_w165, c0_n10_w166, c0_n10_w167, c0_n10_w168, c0_n10_w169, c0_n10_w170, c0_n10_w171, c0_n10_w172, c0_n10_w173, c0_n10_w174, c0_n10_w175, c0_n10_w176, c0_n10_w177, c0_n10_w178, c0_n10_w179, c0_n10_w180, c0_n10_w181, c0_n10_w182, c0_n10_w183, c0_n10_w184, c0_n10_w185, c0_n10_w186, c0_n10_w187, c0_n10_w188, c0_n10_w189, c0_n10_w190, c0_n10_w191, c0_n10_w192, c0_n10_w193, c0_n10_w194, c0_n10_w195, c0_n10_w196, c0_n10_w197, c0_n10_w198, c0_n10_w199, c0_n10_w200, c0_n11_w1, c0_n11_w2, c0_n11_w3, c0_n11_w4, c0_n11_w5, c0_n11_w6, c0_n11_w7, c0_n11_w8, c0_n11_w9, c0_n11_w10, c0_n11_w11, c0_n11_w12, c0_n11_w13, c0_n11_w14, c0_n11_w15, c0_n11_w16, c0_n11_w17, c0_n11_w18, c0_n11_w19, c0_n11_w20, c0_n11_w21, c0_n11_w22, c0_n11_w23, c0_n11_w24, c0_n11_w25, c0_n11_w26, c0_n11_w27, c0_n11_w28, c0_n11_w29, c0_n11_w30, c0_n11_w31, c0_n11_w32, c0_n11_w33, c0_n11_w34, c0_n11_w35, c0_n11_w36, c0_n11_w37, c0_n11_w38, c0_n11_w39, c0_n11_w40, c0_n11_w41, c0_n11_w42, c0_n11_w43, c0_n11_w44, c0_n11_w45, c0_n11_w46, c0_n11_w47, c0_n11_w48, c0_n11_w49, c0_n11_w50, c0_n11_w51, c0_n11_w52, c0_n11_w53, c0_n11_w54, c0_n11_w55, c0_n11_w56, c0_n11_w57, c0_n11_w58, c0_n11_w59, c0_n11_w60, c0_n11_w61, c0_n11_w62, c0_n11_w63, c0_n11_w64, c0_n11_w65, c0_n11_w66, c0_n11_w67, c0_n11_w68, c0_n11_w69, c0_n11_w70, c0_n11_w71, c0_n11_w72, c0_n11_w73, c0_n11_w74, c0_n11_w75, c0_n11_w76, c0_n11_w77, c0_n11_w78, c0_n11_w79, c0_n11_w80, c0_n11_w81, c0_n11_w82, c0_n11_w83, c0_n11_w84, c0_n11_w85, c0_n11_w86, c0_n11_w87, c0_n11_w88, c0_n11_w89, c0_n11_w90, c0_n11_w91, c0_n11_w92, c0_n11_w93, c0_n11_w94, c0_n11_w95, c0_n11_w96, c0_n11_w97, c0_n11_w98, c0_n11_w99, c0_n11_w100, c0_n11_w101, c0_n11_w102, c0_n11_w103, c0_n11_w104, c0_n11_w105, c0_n11_w106, c0_n11_w107, c0_n11_w108, c0_n11_w109, c0_n11_w110, c0_n11_w111, c0_n11_w112, c0_n11_w113, c0_n11_w114, c0_n11_w115, c0_n11_w116, c0_n11_w117, c0_n11_w118, c0_n11_w119, c0_n11_w120, c0_n11_w121, c0_n11_w122, c0_n11_w123, c0_n11_w124, c0_n11_w125, c0_n11_w126, c0_n11_w127, c0_n11_w128, c0_n11_w129, c0_n11_w130, c0_n11_w131, c0_n11_w132, c0_n11_w133, c0_n11_w134, c0_n11_w135, c0_n11_w136, c0_n11_w137, c0_n11_w138, c0_n11_w139, c0_n11_w140, c0_n11_w141, c0_n11_w142, c0_n11_w143, c0_n11_w144, c0_n11_w145, c0_n11_w146, c0_n11_w147, c0_n11_w148, c0_n11_w149, c0_n11_w150, c0_n11_w151, c0_n11_w152, c0_n11_w153, c0_n11_w154, c0_n11_w155, c0_n11_w156, c0_n11_w157, c0_n11_w158, c0_n11_w159, c0_n11_w160, c0_n11_w161, c0_n11_w162, c0_n11_w163, c0_n11_w164, c0_n11_w165, c0_n11_w166, c0_n11_w167, c0_n11_w168, c0_n11_w169, c0_n11_w170, c0_n11_w171, c0_n11_w172, c0_n11_w173, c0_n11_w174, c0_n11_w175, c0_n11_w176, c0_n11_w177, c0_n11_w178, c0_n11_w179, c0_n11_w180, c0_n11_w181, c0_n11_w182, c0_n11_w183, c0_n11_w184, c0_n11_w185, c0_n11_w186, c0_n11_w187, c0_n11_w188, c0_n11_w189, c0_n11_w190, c0_n11_w191, c0_n11_w192, c0_n11_w193, c0_n11_w194, c0_n11_w195, c0_n11_w196, c0_n11_w197, c0_n11_w198, c0_n11_w199, c0_n11_w200, c0_n12_w1, c0_n12_w2, c0_n12_w3, c0_n12_w4, c0_n12_w5, c0_n12_w6, c0_n12_w7, c0_n12_w8, c0_n12_w9, c0_n12_w10, c0_n12_w11, c0_n12_w12, c0_n12_w13, c0_n12_w14, c0_n12_w15, c0_n12_w16, c0_n12_w17, c0_n12_w18, c0_n12_w19, c0_n12_w20, c0_n12_w21, c0_n12_w22, c0_n12_w23, c0_n12_w24, c0_n12_w25, c0_n12_w26, c0_n12_w27, c0_n12_w28, c0_n12_w29, c0_n12_w30, c0_n12_w31, c0_n12_w32, c0_n12_w33, c0_n12_w34, c0_n12_w35, c0_n12_w36, c0_n12_w37, c0_n12_w38, c0_n12_w39, c0_n12_w40, c0_n12_w41, c0_n12_w42, c0_n12_w43, c0_n12_w44, c0_n12_w45, c0_n12_w46, c0_n12_w47, c0_n12_w48, c0_n12_w49, c0_n12_w50, c0_n12_w51, c0_n12_w52, c0_n12_w53, c0_n12_w54, c0_n12_w55, c0_n12_w56, c0_n12_w57, c0_n12_w58, c0_n12_w59, c0_n12_w60, c0_n12_w61, c0_n12_w62, c0_n12_w63, c0_n12_w64, c0_n12_w65, c0_n12_w66, c0_n12_w67, c0_n12_w68, c0_n12_w69, c0_n12_w70, c0_n12_w71, c0_n12_w72, c0_n12_w73, c0_n12_w74, c0_n12_w75, c0_n12_w76, c0_n12_w77, c0_n12_w78, c0_n12_w79, c0_n12_w80, c0_n12_w81, c0_n12_w82, c0_n12_w83, c0_n12_w84, c0_n12_w85, c0_n12_w86, c0_n12_w87, c0_n12_w88, c0_n12_w89, c0_n12_w90, c0_n12_w91, c0_n12_w92, c0_n12_w93, c0_n12_w94, c0_n12_w95, c0_n12_w96, c0_n12_w97, c0_n12_w98, c0_n12_w99, c0_n12_w100, c0_n12_w101, c0_n12_w102, c0_n12_w103, c0_n12_w104, c0_n12_w105, c0_n12_w106, c0_n12_w107, c0_n12_w108, c0_n12_w109, c0_n12_w110, c0_n12_w111, c0_n12_w112, c0_n12_w113, c0_n12_w114, c0_n12_w115, c0_n12_w116, c0_n12_w117, c0_n12_w118, c0_n12_w119, c0_n12_w120, c0_n12_w121, c0_n12_w122, c0_n12_w123, c0_n12_w124, c0_n12_w125, c0_n12_w126, c0_n12_w127, c0_n12_w128, c0_n12_w129, c0_n12_w130, c0_n12_w131, c0_n12_w132, c0_n12_w133, c0_n12_w134, c0_n12_w135, c0_n12_w136, c0_n12_w137, c0_n12_w138, c0_n12_w139, c0_n12_w140, c0_n12_w141, c0_n12_w142, c0_n12_w143, c0_n12_w144, c0_n12_w145, c0_n12_w146, c0_n12_w147, c0_n12_w148, c0_n12_w149, c0_n12_w150, c0_n12_w151, c0_n12_w152, c0_n12_w153, c0_n12_w154, c0_n12_w155, c0_n12_w156, c0_n12_w157, c0_n12_w158, c0_n12_w159, c0_n12_w160, c0_n12_w161, c0_n12_w162, c0_n12_w163, c0_n12_w164, c0_n12_w165, c0_n12_w166, c0_n12_w167, c0_n12_w168, c0_n12_w169, c0_n12_w170, c0_n12_w171, c0_n12_w172, c0_n12_w173, c0_n12_w174, c0_n12_w175, c0_n12_w176, c0_n12_w177, c0_n12_w178, c0_n12_w179, c0_n12_w180, c0_n12_w181, c0_n12_w182, c0_n12_w183, c0_n12_w184, c0_n12_w185, c0_n12_w186, c0_n12_w187, c0_n12_w188, c0_n12_w189, c0_n12_w190, c0_n12_w191, c0_n12_w192, c0_n12_w193, c0_n12_w194, c0_n12_w195, c0_n12_w196, c0_n12_w197, c0_n12_w198, c0_n12_w199, c0_n12_w200, c0_n13_w1, c0_n13_w2, c0_n13_w3, c0_n13_w4, c0_n13_w5, c0_n13_w6, c0_n13_w7, c0_n13_w8, c0_n13_w9, c0_n13_w10, c0_n13_w11, c0_n13_w12, c0_n13_w13, c0_n13_w14, c0_n13_w15, c0_n13_w16, c0_n13_w17, c0_n13_w18, c0_n13_w19, c0_n13_w20, c0_n13_w21, c0_n13_w22, c0_n13_w23, c0_n13_w24, c0_n13_w25, c0_n13_w26, c0_n13_w27, c0_n13_w28, c0_n13_w29, c0_n13_w30, c0_n13_w31, c0_n13_w32, c0_n13_w33, c0_n13_w34, c0_n13_w35, c0_n13_w36, c0_n13_w37, c0_n13_w38, c0_n13_w39, c0_n13_w40, c0_n13_w41, c0_n13_w42, c0_n13_w43, c0_n13_w44, c0_n13_w45, c0_n13_w46, c0_n13_w47, c0_n13_w48, c0_n13_w49, c0_n13_w50, c0_n13_w51, c0_n13_w52, c0_n13_w53, c0_n13_w54, c0_n13_w55, c0_n13_w56, c0_n13_w57, c0_n13_w58, c0_n13_w59, c0_n13_w60, c0_n13_w61, c0_n13_w62, c0_n13_w63, c0_n13_w64, c0_n13_w65, c0_n13_w66, c0_n13_w67, c0_n13_w68, c0_n13_w69, c0_n13_w70, c0_n13_w71, c0_n13_w72, c0_n13_w73, c0_n13_w74, c0_n13_w75, c0_n13_w76, c0_n13_w77, c0_n13_w78, c0_n13_w79, c0_n13_w80, c0_n13_w81, c0_n13_w82, c0_n13_w83, c0_n13_w84, c0_n13_w85, c0_n13_w86, c0_n13_w87, c0_n13_w88, c0_n13_w89, c0_n13_w90, c0_n13_w91, c0_n13_w92, c0_n13_w93, c0_n13_w94, c0_n13_w95, c0_n13_w96, c0_n13_w97, c0_n13_w98, c0_n13_w99, c0_n13_w100, c0_n13_w101, c0_n13_w102, c0_n13_w103, c0_n13_w104, c0_n13_w105, c0_n13_w106, c0_n13_w107, c0_n13_w108, c0_n13_w109, c0_n13_w110, c0_n13_w111, c0_n13_w112, c0_n13_w113, c0_n13_w114, c0_n13_w115, c0_n13_w116, c0_n13_w117, c0_n13_w118, c0_n13_w119, c0_n13_w120, c0_n13_w121, c0_n13_w122, c0_n13_w123, c0_n13_w124, c0_n13_w125, c0_n13_w126, c0_n13_w127, c0_n13_w128, c0_n13_w129, c0_n13_w130, c0_n13_w131, c0_n13_w132, c0_n13_w133, c0_n13_w134, c0_n13_w135, c0_n13_w136, c0_n13_w137, c0_n13_w138, c0_n13_w139, c0_n13_w140, c0_n13_w141, c0_n13_w142, c0_n13_w143, c0_n13_w144, c0_n13_w145, c0_n13_w146, c0_n13_w147, c0_n13_w148, c0_n13_w149, c0_n13_w150, c0_n13_w151, c0_n13_w152, c0_n13_w153, c0_n13_w154, c0_n13_w155, c0_n13_w156, c0_n13_w157, c0_n13_w158, c0_n13_w159, c0_n13_w160, c0_n13_w161, c0_n13_w162, c0_n13_w163, c0_n13_w164, c0_n13_w165, c0_n13_w166, c0_n13_w167, c0_n13_w168, c0_n13_w169, c0_n13_w170, c0_n13_w171, c0_n13_w172, c0_n13_w173, c0_n13_w174, c0_n13_w175, c0_n13_w176, c0_n13_w177, c0_n13_w178, c0_n13_w179, c0_n13_w180, c0_n13_w181, c0_n13_w182, c0_n13_w183, c0_n13_w184, c0_n13_w185, c0_n13_w186, c0_n13_w187, c0_n13_w188, c0_n13_w189, c0_n13_w190, c0_n13_w191, c0_n13_w192, c0_n13_w193, c0_n13_w194, c0_n13_w195, c0_n13_w196, c0_n13_w197, c0_n13_w198, c0_n13_w199, c0_n13_w200, c0_n14_w1, c0_n14_w2, c0_n14_w3, c0_n14_w4, c0_n14_w5, c0_n14_w6, c0_n14_w7, c0_n14_w8, c0_n14_w9, c0_n14_w10, c0_n14_w11, c0_n14_w12, c0_n14_w13, c0_n14_w14, c0_n14_w15, c0_n14_w16, c0_n14_w17, c0_n14_w18, c0_n14_w19, c0_n14_w20, c0_n14_w21, c0_n14_w22, c0_n14_w23, c0_n14_w24, c0_n14_w25, c0_n14_w26, c0_n14_w27, c0_n14_w28, c0_n14_w29, c0_n14_w30, c0_n14_w31, c0_n14_w32, c0_n14_w33, c0_n14_w34, c0_n14_w35, c0_n14_w36, c0_n14_w37, c0_n14_w38, c0_n14_w39, c0_n14_w40, c0_n14_w41, c0_n14_w42, c0_n14_w43, c0_n14_w44, c0_n14_w45, c0_n14_w46, c0_n14_w47, c0_n14_w48, c0_n14_w49, c0_n14_w50, c0_n14_w51, c0_n14_w52, c0_n14_w53, c0_n14_w54, c0_n14_w55, c0_n14_w56, c0_n14_w57, c0_n14_w58, c0_n14_w59, c0_n14_w60, c0_n14_w61, c0_n14_w62, c0_n14_w63, c0_n14_w64, c0_n14_w65, c0_n14_w66, c0_n14_w67, c0_n14_w68, c0_n14_w69, c0_n14_w70, c0_n14_w71, c0_n14_w72, c0_n14_w73, c0_n14_w74, c0_n14_w75, c0_n14_w76, c0_n14_w77, c0_n14_w78, c0_n14_w79, c0_n14_w80, c0_n14_w81, c0_n14_w82, c0_n14_w83, c0_n14_w84, c0_n14_w85, c0_n14_w86, c0_n14_w87, c0_n14_w88, c0_n14_w89, c0_n14_w90, c0_n14_w91, c0_n14_w92, c0_n14_w93, c0_n14_w94, c0_n14_w95, c0_n14_w96, c0_n14_w97, c0_n14_w98, c0_n14_w99, c0_n14_w100, c0_n14_w101, c0_n14_w102, c0_n14_w103, c0_n14_w104, c0_n14_w105, c0_n14_w106, c0_n14_w107, c0_n14_w108, c0_n14_w109, c0_n14_w110, c0_n14_w111, c0_n14_w112, c0_n14_w113, c0_n14_w114, c0_n14_w115, c0_n14_w116, c0_n14_w117, c0_n14_w118, c0_n14_w119, c0_n14_w120, c0_n14_w121, c0_n14_w122, c0_n14_w123, c0_n14_w124, c0_n14_w125, c0_n14_w126, c0_n14_w127, c0_n14_w128, c0_n14_w129, c0_n14_w130, c0_n14_w131, c0_n14_w132, c0_n14_w133, c0_n14_w134, c0_n14_w135, c0_n14_w136, c0_n14_w137, c0_n14_w138, c0_n14_w139, c0_n14_w140, c0_n14_w141, c0_n14_w142, c0_n14_w143, c0_n14_w144, c0_n14_w145, c0_n14_w146, c0_n14_w147, c0_n14_w148, c0_n14_w149, c0_n14_w150, c0_n14_w151, c0_n14_w152, c0_n14_w153, c0_n14_w154, c0_n14_w155, c0_n14_w156, c0_n14_w157, c0_n14_w158, c0_n14_w159, c0_n14_w160, c0_n14_w161, c0_n14_w162, c0_n14_w163, c0_n14_w164, c0_n14_w165, c0_n14_w166, c0_n14_w167, c0_n14_w168, c0_n14_w169, c0_n14_w170, c0_n14_w171, c0_n14_w172, c0_n14_w173, c0_n14_w174, c0_n14_w175, c0_n14_w176, c0_n14_w177, c0_n14_w178, c0_n14_w179, c0_n14_w180, c0_n14_w181, c0_n14_w182, c0_n14_w183, c0_n14_w184, c0_n14_w185, c0_n14_w186, c0_n14_w187, c0_n14_w188, c0_n14_w189, c0_n14_w190, c0_n14_w191, c0_n14_w192, c0_n14_w193, c0_n14_w194, c0_n14_w195, c0_n14_w196, c0_n14_w197, c0_n14_w198, c0_n14_w199, c0_n14_w200, c0_n15_w1, c0_n15_w2, c0_n15_w3, c0_n15_w4, c0_n15_w5, c0_n15_w6, c0_n15_w7, c0_n15_w8, c0_n15_w9, c0_n15_w10, c0_n15_w11, c0_n15_w12, c0_n15_w13, c0_n15_w14, c0_n15_w15, c0_n15_w16, c0_n15_w17, c0_n15_w18, c0_n15_w19, c0_n15_w20, c0_n15_w21, c0_n15_w22, c0_n15_w23, c0_n15_w24, c0_n15_w25, c0_n15_w26, c0_n15_w27, c0_n15_w28, c0_n15_w29, c0_n15_w30, c0_n15_w31, c0_n15_w32, c0_n15_w33, c0_n15_w34, c0_n15_w35, c0_n15_w36, c0_n15_w37, c0_n15_w38, c0_n15_w39, c0_n15_w40, c0_n15_w41, c0_n15_w42, c0_n15_w43, c0_n15_w44, c0_n15_w45, c0_n15_w46, c0_n15_w47, c0_n15_w48, c0_n15_w49, c0_n15_w50, c0_n15_w51, c0_n15_w52, c0_n15_w53, c0_n15_w54, c0_n15_w55, c0_n15_w56, c0_n15_w57, c0_n15_w58, c0_n15_w59, c0_n15_w60, c0_n15_w61, c0_n15_w62, c0_n15_w63, c0_n15_w64, c0_n15_w65, c0_n15_w66, c0_n15_w67, c0_n15_w68, c0_n15_w69, c0_n15_w70, c0_n15_w71, c0_n15_w72, c0_n15_w73, c0_n15_w74, c0_n15_w75, c0_n15_w76, c0_n15_w77, c0_n15_w78, c0_n15_w79, c0_n15_w80, c0_n15_w81, c0_n15_w82, c0_n15_w83, c0_n15_w84, c0_n15_w85, c0_n15_w86, c0_n15_w87, c0_n15_w88, c0_n15_w89, c0_n15_w90, c0_n15_w91, c0_n15_w92, c0_n15_w93, c0_n15_w94, c0_n15_w95, c0_n15_w96, c0_n15_w97, c0_n15_w98, c0_n15_w99, c0_n15_w100, c0_n15_w101, c0_n15_w102, c0_n15_w103, c0_n15_w104, c0_n15_w105, c0_n15_w106, c0_n15_w107, c0_n15_w108, c0_n15_w109, c0_n15_w110, c0_n15_w111, c0_n15_w112, c0_n15_w113, c0_n15_w114, c0_n15_w115, c0_n15_w116, c0_n15_w117, c0_n15_w118, c0_n15_w119, c0_n15_w120, c0_n15_w121, c0_n15_w122, c0_n15_w123, c0_n15_w124, c0_n15_w125, c0_n15_w126, c0_n15_w127, c0_n15_w128, c0_n15_w129, c0_n15_w130, c0_n15_w131, c0_n15_w132, c0_n15_w133, c0_n15_w134, c0_n15_w135, c0_n15_w136, c0_n15_w137, c0_n15_w138, c0_n15_w139, c0_n15_w140, c0_n15_w141, c0_n15_w142, c0_n15_w143, c0_n15_w144, c0_n15_w145, c0_n15_w146, c0_n15_w147, c0_n15_w148, c0_n15_w149, c0_n15_w150, c0_n15_w151, c0_n15_w152, c0_n15_w153, c0_n15_w154, c0_n15_w155, c0_n15_w156, c0_n15_w157, c0_n15_w158, c0_n15_w159, c0_n15_w160, c0_n15_w161, c0_n15_w162, c0_n15_w163, c0_n15_w164, c0_n15_w165, c0_n15_w166, c0_n15_w167, c0_n15_w168, c0_n15_w169, c0_n15_w170, c0_n15_w171, c0_n15_w172, c0_n15_w173, c0_n15_w174, c0_n15_w175, c0_n15_w176, c0_n15_w177, c0_n15_w178, c0_n15_w179, c0_n15_w180, c0_n15_w181, c0_n15_w182, c0_n15_w183, c0_n15_w184, c0_n15_w185, c0_n15_w186, c0_n15_w187, c0_n15_w188, c0_n15_w189, c0_n15_w190, c0_n15_w191, c0_n15_w192, c0_n15_w193, c0_n15_w194, c0_n15_w195, c0_n15_w196, c0_n15_w197, c0_n15_w198, c0_n15_w199, c0_n15_w200, c0_n16_w1, c0_n16_w2, c0_n16_w3, c0_n16_w4, c0_n16_w5, c0_n16_w6, c0_n16_w7, c0_n16_w8, c0_n16_w9, c0_n16_w10, c0_n16_w11, c0_n16_w12, c0_n16_w13, c0_n16_w14, c0_n16_w15, c0_n16_w16, c0_n16_w17, c0_n16_w18, c0_n16_w19, c0_n16_w20, c0_n16_w21, c0_n16_w22, c0_n16_w23, c0_n16_w24, c0_n16_w25, c0_n16_w26, c0_n16_w27, c0_n16_w28, c0_n16_w29, c0_n16_w30, c0_n16_w31, c0_n16_w32, c0_n16_w33, c0_n16_w34, c0_n16_w35, c0_n16_w36, c0_n16_w37, c0_n16_w38, c0_n16_w39, c0_n16_w40, c0_n16_w41, c0_n16_w42, c0_n16_w43, c0_n16_w44, c0_n16_w45, c0_n16_w46, c0_n16_w47, c0_n16_w48, c0_n16_w49, c0_n16_w50, c0_n16_w51, c0_n16_w52, c0_n16_w53, c0_n16_w54, c0_n16_w55, c0_n16_w56, c0_n16_w57, c0_n16_w58, c0_n16_w59, c0_n16_w60, c0_n16_w61, c0_n16_w62, c0_n16_w63, c0_n16_w64, c0_n16_w65, c0_n16_w66, c0_n16_w67, c0_n16_w68, c0_n16_w69, c0_n16_w70, c0_n16_w71, c0_n16_w72, c0_n16_w73, c0_n16_w74, c0_n16_w75, c0_n16_w76, c0_n16_w77, c0_n16_w78, c0_n16_w79, c0_n16_w80, c0_n16_w81, c0_n16_w82, c0_n16_w83, c0_n16_w84, c0_n16_w85, c0_n16_w86, c0_n16_w87, c0_n16_w88, c0_n16_w89, c0_n16_w90, c0_n16_w91, c0_n16_w92, c0_n16_w93, c0_n16_w94, c0_n16_w95, c0_n16_w96, c0_n16_w97, c0_n16_w98, c0_n16_w99, c0_n16_w100, c0_n16_w101, c0_n16_w102, c0_n16_w103, c0_n16_w104, c0_n16_w105, c0_n16_w106, c0_n16_w107, c0_n16_w108, c0_n16_w109, c0_n16_w110, c0_n16_w111, c0_n16_w112, c0_n16_w113, c0_n16_w114, c0_n16_w115, c0_n16_w116, c0_n16_w117, c0_n16_w118, c0_n16_w119, c0_n16_w120, c0_n16_w121, c0_n16_w122, c0_n16_w123, c0_n16_w124, c0_n16_w125, c0_n16_w126, c0_n16_w127, c0_n16_w128, c0_n16_w129, c0_n16_w130, c0_n16_w131, c0_n16_w132, c0_n16_w133, c0_n16_w134, c0_n16_w135, c0_n16_w136, c0_n16_w137, c0_n16_w138, c0_n16_w139, c0_n16_w140, c0_n16_w141, c0_n16_w142, c0_n16_w143, c0_n16_w144, c0_n16_w145, c0_n16_w146, c0_n16_w147, c0_n16_w148, c0_n16_w149, c0_n16_w150, c0_n16_w151, c0_n16_w152, c0_n16_w153, c0_n16_w154, c0_n16_w155, c0_n16_w156, c0_n16_w157, c0_n16_w158, c0_n16_w159, c0_n16_w160, c0_n16_w161, c0_n16_w162, c0_n16_w163, c0_n16_w164, c0_n16_w165, c0_n16_w166, c0_n16_w167, c0_n16_w168, c0_n16_w169, c0_n16_w170, c0_n16_w171, c0_n16_w172, c0_n16_w173, c0_n16_w174, c0_n16_w175, c0_n16_w176, c0_n16_w177, c0_n16_w178, c0_n16_w179, c0_n16_w180, c0_n16_w181, c0_n16_w182, c0_n16_w183, c0_n16_w184, c0_n16_w185, c0_n16_w186, c0_n16_w187, c0_n16_w188, c0_n16_w189, c0_n16_w190, c0_n16_w191, c0_n16_w192, c0_n16_w193, c0_n16_w194, c0_n16_w195, c0_n16_w196, c0_n16_w197, c0_n16_w198, c0_n16_w199, c0_n16_w200, c0_n17_w1, c0_n17_w2, c0_n17_w3, c0_n17_w4, c0_n17_w5, c0_n17_w6, c0_n17_w7, c0_n17_w8, c0_n17_w9, c0_n17_w10, c0_n17_w11, c0_n17_w12, c0_n17_w13, c0_n17_w14, c0_n17_w15, c0_n17_w16, c0_n17_w17, c0_n17_w18, c0_n17_w19, c0_n17_w20, c0_n17_w21, c0_n17_w22, c0_n17_w23, c0_n17_w24, c0_n17_w25, c0_n17_w26, c0_n17_w27, c0_n17_w28, c0_n17_w29, c0_n17_w30, c0_n17_w31, c0_n17_w32, c0_n17_w33, c0_n17_w34, c0_n17_w35, c0_n17_w36, c0_n17_w37, c0_n17_w38, c0_n17_w39, c0_n17_w40, c0_n17_w41, c0_n17_w42, c0_n17_w43, c0_n17_w44, c0_n17_w45, c0_n17_w46, c0_n17_w47, c0_n17_w48, c0_n17_w49, c0_n17_w50, c0_n17_w51, c0_n17_w52, c0_n17_w53, c0_n17_w54, c0_n17_w55, c0_n17_w56, c0_n17_w57, c0_n17_w58, c0_n17_w59, c0_n17_w60, c0_n17_w61, c0_n17_w62, c0_n17_w63, c0_n17_w64, c0_n17_w65, c0_n17_w66, c0_n17_w67, c0_n17_w68, c0_n17_w69, c0_n17_w70, c0_n17_w71, c0_n17_w72, c0_n17_w73, c0_n17_w74, c0_n17_w75, c0_n17_w76, c0_n17_w77, c0_n17_w78, c0_n17_w79, c0_n17_w80, c0_n17_w81, c0_n17_w82, c0_n17_w83, c0_n17_w84, c0_n17_w85, c0_n17_w86, c0_n17_w87, c0_n17_w88, c0_n17_w89, c0_n17_w90, c0_n17_w91, c0_n17_w92, c0_n17_w93, c0_n17_w94, c0_n17_w95, c0_n17_w96, c0_n17_w97, c0_n17_w98, c0_n17_w99, c0_n17_w100, c0_n17_w101, c0_n17_w102, c0_n17_w103, c0_n17_w104, c0_n17_w105, c0_n17_w106, c0_n17_w107, c0_n17_w108, c0_n17_w109, c0_n17_w110, c0_n17_w111, c0_n17_w112, c0_n17_w113, c0_n17_w114, c0_n17_w115, c0_n17_w116, c0_n17_w117, c0_n17_w118, c0_n17_w119, c0_n17_w120, c0_n17_w121, c0_n17_w122, c0_n17_w123, c0_n17_w124, c0_n17_w125, c0_n17_w126, c0_n17_w127, c0_n17_w128, c0_n17_w129, c0_n17_w130, c0_n17_w131, c0_n17_w132, c0_n17_w133, c0_n17_w134, c0_n17_w135, c0_n17_w136, c0_n17_w137, c0_n17_w138, c0_n17_w139, c0_n17_w140, c0_n17_w141, c0_n17_w142, c0_n17_w143, c0_n17_w144, c0_n17_w145, c0_n17_w146, c0_n17_w147, c0_n17_w148, c0_n17_w149, c0_n17_w150, c0_n17_w151, c0_n17_w152, c0_n17_w153, c0_n17_w154, c0_n17_w155, c0_n17_w156, c0_n17_w157, c0_n17_w158, c0_n17_w159, c0_n17_w160, c0_n17_w161, c0_n17_w162, c0_n17_w163, c0_n17_w164, c0_n17_w165, c0_n17_w166, c0_n17_w167, c0_n17_w168, c0_n17_w169, c0_n17_w170, c0_n17_w171, c0_n17_w172, c0_n17_w173, c0_n17_w174, c0_n17_w175, c0_n17_w176, c0_n17_w177, c0_n17_w178, c0_n17_w179, c0_n17_w180, c0_n17_w181, c0_n17_w182, c0_n17_w183, c0_n17_w184, c0_n17_w185, c0_n17_w186, c0_n17_w187, c0_n17_w188, c0_n17_w189, c0_n17_w190, c0_n17_w191, c0_n17_w192, c0_n17_w193, c0_n17_w194, c0_n17_w195, c0_n17_w196, c0_n17_w197, c0_n17_w198, c0_n17_w199, c0_n17_w200, c0_n18_w1, c0_n18_w2, c0_n18_w3, c0_n18_w4, c0_n18_w5, c0_n18_w6, c0_n18_w7, c0_n18_w8, c0_n18_w9, c0_n18_w10, c0_n18_w11, c0_n18_w12, c0_n18_w13, c0_n18_w14, c0_n18_w15, c0_n18_w16, c0_n18_w17, c0_n18_w18, c0_n18_w19, c0_n18_w20, c0_n18_w21, c0_n18_w22, c0_n18_w23, c0_n18_w24, c0_n18_w25, c0_n18_w26, c0_n18_w27, c0_n18_w28, c0_n18_w29, c0_n18_w30, c0_n18_w31, c0_n18_w32, c0_n18_w33, c0_n18_w34, c0_n18_w35, c0_n18_w36, c0_n18_w37, c0_n18_w38, c0_n18_w39, c0_n18_w40, c0_n18_w41, c0_n18_w42, c0_n18_w43, c0_n18_w44, c0_n18_w45, c0_n18_w46, c0_n18_w47, c0_n18_w48, c0_n18_w49, c0_n18_w50, c0_n18_w51, c0_n18_w52, c0_n18_w53, c0_n18_w54, c0_n18_w55, c0_n18_w56, c0_n18_w57, c0_n18_w58, c0_n18_w59, c0_n18_w60, c0_n18_w61, c0_n18_w62, c0_n18_w63, c0_n18_w64, c0_n18_w65, c0_n18_w66, c0_n18_w67, c0_n18_w68, c0_n18_w69, c0_n18_w70, c0_n18_w71, c0_n18_w72, c0_n18_w73, c0_n18_w74, c0_n18_w75, c0_n18_w76, c0_n18_w77, c0_n18_w78, c0_n18_w79, c0_n18_w80, c0_n18_w81, c0_n18_w82, c0_n18_w83, c0_n18_w84, c0_n18_w85, c0_n18_w86, c0_n18_w87, c0_n18_w88, c0_n18_w89, c0_n18_w90, c0_n18_w91, c0_n18_w92, c0_n18_w93, c0_n18_w94, c0_n18_w95, c0_n18_w96, c0_n18_w97, c0_n18_w98, c0_n18_w99, c0_n18_w100, c0_n18_w101, c0_n18_w102, c0_n18_w103, c0_n18_w104, c0_n18_w105, c0_n18_w106, c0_n18_w107, c0_n18_w108, c0_n18_w109, c0_n18_w110, c0_n18_w111, c0_n18_w112, c0_n18_w113, c0_n18_w114, c0_n18_w115, c0_n18_w116, c0_n18_w117, c0_n18_w118, c0_n18_w119, c0_n18_w120, c0_n18_w121, c0_n18_w122, c0_n18_w123, c0_n18_w124, c0_n18_w125, c0_n18_w126, c0_n18_w127, c0_n18_w128, c0_n18_w129, c0_n18_w130, c0_n18_w131, c0_n18_w132, c0_n18_w133, c0_n18_w134, c0_n18_w135, c0_n18_w136, c0_n18_w137, c0_n18_w138, c0_n18_w139, c0_n18_w140, c0_n18_w141, c0_n18_w142, c0_n18_w143, c0_n18_w144, c0_n18_w145, c0_n18_w146, c0_n18_w147, c0_n18_w148, c0_n18_w149, c0_n18_w150, c0_n18_w151, c0_n18_w152, c0_n18_w153, c0_n18_w154, c0_n18_w155, c0_n18_w156, c0_n18_w157, c0_n18_w158, c0_n18_w159, c0_n18_w160, c0_n18_w161, c0_n18_w162, c0_n18_w163, c0_n18_w164, c0_n18_w165, c0_n18_w166, c0_n18_w167, c0_n18_w168, c0_n18_w169, c0_n18_w170, c0_n18_w171, c0_n18_w172, c0_n18_w173, c0_n18_w174, c0_n18_w175, c0_n18_w176, c0_n18_w177, c0_n18_w178, c0_n18_w179, c0_n18_w180, c0_n18_w181, c0_n18_w182, c0_n18_w183, c0_n18_w184, c0_n18_w185, c0_n18_w186, c0_n18_w187, c0_n18_w188, c0_n18_w189, c0_n18_w190, c0_n18_w191, c0_n18_w192, c0_n18_w193, c0_n18_w194, c0_n18_w195, c0_n18_w196, c0_n18_w197, c0_n18_w198, c0_n18_w199, c0_n18_w200, c0_n19_w1, c0_n19_w2, c0_n19_w3, c0_n19_w4, c0_n19_w5, c0_n19_w6, c0_n19_w7, c0_n19_w8, c0_n19_w9, c0_n19_w10, c0_n19_w11, c0_n19_w12, c0_n19_w13, c0_n19_w14, c0_n19_w15, c0_n19_w16, c0_n19_w17, c0_n19_w18, c0_n19_w19, c0_n19_w20, c0_n19_w21, c0_n19_w22, c0_n19_w23, c0_n19_w24, c0_n19_w25, c0_n19_w26, c0_n19_w27, c0_n19_w28, c0_n19_w29, c0_n19_w30, c0_n19_w31, c0_n19_w32, c0_n19_w33, c0_n19_w34, c0_n19_w35, c0_n19_w36, c0_n19_w37, c0_n19_w38, c0_n19_w39, c0_n19_w40, c0_n19_w41, c0_n19_w42, c0_n19_w43, c0_n19_w44, c0_n19_w45, c0_n19_w46, c0_n19_w47, c0_n19_w48, c0_n19_w49, c0_n19_w50, c0_n19_w51, c0_n19_w52, c0_n19_w53, c0_n19_w54, c0_n19_w55, c0_n19_w56, c0_n19_w57, c0_n19_w58, c0_n19_w59, c0_n19_w60, c0_n19_w61, c0_n19_w62, c0_n19_w63, c0_n19_w64, c0_n19_w65, c0_n19_w66, c0_n19_w67, c0_n19_w68, c0_n19_w69, c0_n19_w70, c0_n19_w71, c0_n19_w72, c0_n19_w73, c0_n19_w74, c0_n19_w75, c0_n19_w76, c0_n19_w77, c0_n19_w78, c0_n19_w79, c0_n19_w80, c0_n19_w81, c0_n19_w82, c0_n19_w83, c0_n19_w84, c0_n19_w85, c0_n19_w86, c0_n19_w87, c0_n19_w88, c0_n19_w89, c0_n19_w90, c0_n19_w91, c0_n19_w92, c0_n19_w93, c0_n19_w94, c0_n19_w95, c0_n19_w96, c0_n19_w97, c0_n19_w98, c0_n19_w99, c0_n19_w100, c0_n19_w101, c0_n19_w102, c0_n19_w103, c0_n19_w104, c0_n19_w105, c0_n19_w106, c0_n19_w107, c0_n19_w108, c0_n19_w109, c0_n19_w110, c0_n19_w111, c0_n19_w112, c0_n19_w113, c0_n19_w114, c0_n19_w115, c0_n19_w116, c0_n19_w117, c0_n19_w118, c0_n19_w119, c0_n19_w120, c0_n19_w121, c0_n19_w122, c0_n19_w123, c0_n19_w124, c0_n19_w125, c0_n19_w126, c0_n19_w127, c0_n19_w128, c0_n19_w129, c0_n19_w130, c0_n19_w131, c0_n19_w132, c0_n19_w133, c0_n19_w134, c0_n19_w135, c0_n19_w136, c0_n19_w137, c0_n19_w138, c0_n19_w139, c0_n19_w140, c0_n19_w141, c0_n19_w142, c0_n19_w143, c0_n19_w144, c0_n19_w145, c0_n19_w146, c0_n19_w147, c0_n19_w148, c0_n19_w149, c0_n19_w150, c0_n19_w151, c0_n19_w152, c0_n19_w153, c0_n19_w154, c0_n19_w155, c0_n19_w156, c0_n19_w157, c0_n19_w158, c0_n19_w159, c0_n19_w160, c0_n19_w161, c0_n19_w162, c0_n19_w163, c0_n19_w164, c0_n19_w165, c0_n19_w166, c0_n19_w167, c0_n19_w168, c0_n19_w169, c0_n19_w170, c0_n19_w171, c0_n19_w172, c0_n19_w173, c0_n19_w174, c0_n19_w175, c0_n19_w176, c0_n19_w177, c0_n19_w178, c0_n19_w179, c0_n19_w180, c0_n19_w181, c0_n19_w182, c0_n19_w183, c0_n19_w184, c0_n19_w185, c0_n19_w186, c0_n19_w187, c0_n19_w188, c0_n19_w189, c0_n19_w190, c0_n19_w191, c0_n19_w192, c0_n19_w193, c0_n19_w194, c0_n19_w195, c0_n19_w196, c0_n19_w197, c0_n19_w198, c0_n19_w199, c0_n19_w200, c0_n20_w1, c0_n20_w2, c0_n20_w3, c0_n20_w4, c0_n20_w5, c0_n20_w6, c0_n20_w7, c0_n20_w8, c0_n20_w9, c0_n20_w10, c0_n20_w11, c0_n20_w12, c0_n20_w13, c0_n20_w14, c0_n20_w15, c0_n20_w16, c0_n20_w17, c0_n20_w18, c0_n20_w19, c0_n20_w20, c0_n20_w21, c0_n20_w22, c0_n20_w23, c0_n20_w24, c0_n20_w25, c0_n20_w26, c0_n20_w27, c0_n20_w28, c0_n20_w29, c0_n20_w30, c0_n20_w31, c0_n20_w32, c0_n20_w33, c0_n20_w34, c0_n20_w35, c0_n20_w36, c0_n20_w37, c0_n20_w38, c0_n20_w39, c0_n20_w40, c0_n20_w41, c0_n20_w42, c0_n20_w43, c0_n20_w44, c0_n20_w45, c0_n20_w46, c0_n20_w47, c0_n20_w48, c0_n20_w49, c0_n20_w50, c0_n20_w51, c0_n20_w52, c0_n20_w53, c0_n20_w54, c0_n20_w55, c0_n20_w56, c0_n20_w57, c0_n20_w58, c0_n20_w59, c0_n20_w60, c0_n20_w61, c0_n20_w62, c0_n20_w63, c0_n20_w64, c0_n20_w65, c0_n20_w66, c0_n20_w67, c0_n20_w68, c0_n20_w69, c0_n20_w70, c0_n20_w71, c0_n20_w72, c0_n20_w73, c0_n20_w74, c0_n20_w75, c0_n20_w76, c0_n20_w77, c0_n20_w78, c0_n20_w79, c0_n20_w80, c0_n20_w81, c0_n20_w82, c0_n20_w83, c0_n20_w84, c0_n20_w85, c0_n20_w86, c0_n20_w87, c0_n20_w88, c0_n20_w89, c0_n20_w90, c0_n20_w91, c0_n20_w92, c0_n20_w93, c0_n20_w94, c0_n20_w95, c0_n20_w96, c0_n20_w97, c0_n20_w98, c0_n20_w99, c0_n20_w100, c0_n20_w101, c0_n20_w102, c0_n20_w103, c0_n20_w104, c0_n20_w105, c0_n20_w106, c0_n20_w107, c0_n20_w108, c0_n20_w109, c0_n20_w110, c0_n20_w111, c0_n20_w112, c0_n20_w113, c0_n20_w114, c0_n20_w115, c0_n20_w116, c0_n20_w117, c0_n20_w118, c0_n20_w119, c0_n20_w120, c0_n20_w121, c0_n20_w122, c0_n20_w123, c0_n20_w124, c0_n20_w125, c0_n20_w126, c0_n20_w127, c0_n20_w128, c0_n20_w129, c0_n20_w130, c0_n20_w131, c0_n20_w132, c0_n20_w133, c0_n20_w134, c0_n20_w135, c0_n20_w136, c0_n20_w137, c0_n20_w138, c0_n20_w139, c0_n20_w140, c0_n20_w141, c0_n20_w142, c0_n20_w143, c0_n20_w144, c0_n20_w145, c0_n20_w146, c0_n20_w147, c0_n20_w148, c0_n20_w149, c0_n20_w150, c0_n20_w151, c0_n20_w152, c0_n20_w153, c0_n20_w154, c0_n20_w155, c0_n20_w156, c0_n20_w157, c0_n20_w158, c0_n20_w159, c0_n20_w160, c0_n20_w161, c0_n20_w162, c0_n20_w163, c0_n20_w164, c0_n20_w165, c0_n20_w166, c0_n20_w167, c0_n20_w168, c0_n20_w169, c0_n20_w170, c0_n20_w171, c0_n20_w172, c0_n20_w173, c0_n20_w174, c0_n20_w175, c0_n20_w176, c0_n20_w177, c0_n20_w178, c0_n20_w179, c0_n20_w180, c0_n20_w181, c0_n20_w182, c0_n20_w183, c0_n20_w184, c0_n20_w185, c0_n20_w186, c0_n20_w187, c0_n20_w188, c0_n20_w189, c0_n20_w190, c0_n20_w191, c0_n20_w192, c0_n20_w193, c0_n20_w194, c0_n20_w195, c0_n20_w196, c0_n20_w197, c0_n20_w198, c0_n20_w199, c0_n20_w200, c0_n21_w1, c0_n21_w2, c0_n21_w3, c0_n21_w4, c0_n21_w5, c0_n21_w6, c0_n21_w7, c0_n21_w8, c0_n21_w9, c0_n21_w10, c0_n21_w11, c0_n21_w12, c0_n21_w13, c0_n21_w14, c0_n21_w15, c0_n21_w16, c0_n21_w17, c0_n21_w18, c0_n21_w19, c0_n21_w20, c0_n21_w21, c0_n21_w22, c0_n21_w23, c0_n21_w24, c0_n21_w25, c0_n21_w26, c0_n21_w27, c0_n21_w28, c0_n21_w29, c0_n21_w30, c0_n21_w31, c0_n21_w32, c0_n21_w33, c0_n21_w34, c0_n21_w35, c0_n21_w36, c0_n21_w37, c0_n21_w38, c0_n21_w39, c0_n21_w40, c0_n21_w41, c0_n21_w42, c0_n21_w43, c0_n21_w44, c0_n21_w45, c0_n21_w46, c0_n21_w47, c0_n21_w48, c0_n21_w49, c0_n21_w50, c0_n21_w51, c0_n21_w52, c0_n21_w53, c0_n21_w54, c0_n21_w55, c0_n21_w56, c0_n21_w57, c0_n21_w58, c0_n21_w59, c0_n21_w60, c0_n21_w61, c0_n21_w62, c0_n21_w63, c0_n21_w64, c0_n21_w65, c0_n21_w66, c0_n21_w67, c0_n21_w68, c0_n21_w69, c0_n21_w70, c0_n21_w71, c0_n21_w72, c0_n21_w73, c0_n21_w74, c0_n21_w75, c0_n21_w76, c0_n21_w77, c0_n21_w78, c0_n21_w79, c0_n21_w80, c0_n21_w81, c0_n21_w82, c0_n21_w83, c0_n21_w84, c0_n21_w85, c0_n21_w86, c0_n21_w87, c0_n21_w88, c0_n21_w89, c0_n21_w90, c0_n21_w91, c0_n21_w92, c0_n21_w93, c0_n21_w94, c0_n21_w95, c0_n21_w96, c0_n21_w97, c0_n21_w98, c0_n21_w99, c0_n21_w100, c0_n21_w101, c0_n21_w102, c0_n21_w103, c0_n21_w104, c0_n21_w105, c0_n21_w106, c0_n21_w107, c0_n21_w108, c0_n21_w109, c0_n21_w110, c0_n21_w111, c0_n21_w112, c0_n21_w113, c0_n21_w114, c0_n21_w115, c0_n21_w116, c0_n21_w117, c0_n21_w118, c0_n21_w119, c0_n21_w120, c0_n21_w121, c0_n21_w122, c0_n21_w123, c0_n21_w124, c0_n21_w125, c0_n21_w126, c0_n21_w127, c0_n21_w128, c0_n21_w129, c0_n21_w130, c0_n21_w131, c0_n21_w132, c0_n21_w133, c0_n21_w134, c0_n21_w135, c0_n21_w136, c0_n21_w137, c0_n21_w138, c0_n21_w139, c0_n21_w140, c0_n21_w141, c0_n21_w142, c0_n21_w143, c0_n21_w144, c0_n21_w145, c0_n21_w146, c0_n21_w147, c0_n21_w148, c0_n21_w149, c0_n21_w150, c0_n21_w151, c0_n21_w152, c0_n21_w153, c0_n21_w154, c0_n21_w155, c0_n21_w156, c0_n21_w157, c0_n21_w158, c0_n21_w159, c0_n21_w160, c0_n21_w161, c0_n21_w162, c0_n21_w163, c0_n21_w164, c0_n21_w165, c0_n21_w166, c0_n21_w167, c0_n21_w168, c0_n21_w169, c0_n21_w170, c0_n21_w171, c0_n21_w172, c0_n21_w173, c0_n21_w174, c0_n21_w175, c0_n21_w176, c0_n21_w177, c0_n21_w178, c0_n21_w179, c0_n21_w180, c0_n21_w181, c0_n21_w182, c0_n21_w183, c0_n21_w184, c0_n21_w185, c0_n21_w186, c0_n21_w187, c0_n21_w188, c0_n21_w189, c0_n21_w190, c0_n21_w191, c0_n21_w192, c0_n21_w193, c0_n21_w194, c0_n21_w195, c0_n21_w196, c0_n21_w197, c0_n21_w198, c0_n21_w199, c0_n21_w200, c0_n22_w1, c0_n22_w2, c0_n22_w3, c0_n22_w4, c0_n22_w5, c0_n22_w6, c0_n22_w7, c0_n22_w8, c0_n22_w9, c0_n22_w10, c0_n22_w11, c0_n22_w12, c0_n22_w13, c0_n22_w14, c0_n22_w15, c0_n22_w16, c0_n22_w17, c0_n22_w18, c0_n22_w19, c0_n22_w20, c0_n22_w21, c0_n22_w22, c0_n22_w23, c0_n22_w24, c0_n22_w25, c0_n22_w26, c0_n22_w27, c0_n22_w28, c0_n22_w29, c0_n22_w30, c0_n22_w31, c0_n22_w32, c0_n22_w33, c0_n22_w34, c0_n22_w35, c0_n22_w36, c0_n22_w37, c0_n22_w38, c0_n22_w39, c0_n22_w40, c0_n22_w41, c0_n22_w42, c0_n22_w43, c0_n22_w44, c0_n22_w45, c0_n22_w46, c0_n22_w47, c0_n22_w48, c0_n22_w49, c0_n22_w50, c0_n22_w51, c0_n22_w52, c0_n22_w53, c0_n22_w54, c0_n22_w55, c0_n22_w56, c0_n22_w57, c0_n22_w58, c0_n22_w59, c0_n22_w60, c0_n22_w61, c0_n22_w62, c0_n22_w63, c0_n22_w64, c0_n22_w65, c0_n22_w66, c0_n22_w67, c0_n22_w68, c0_n22_w69, c0_n22_w70, c0_n22_w71, c0_n22_w72, c0_n22_w73, c0_n22_w74, c0_n22_w75, c0_n22_w76, c0_n22_w77, c0_n22_w78, c0_n22_w79, c0_n22_w80, c0_n22_w81, c0_n22_w82, c0_n22_w83, c0_n22_w84, c0_n22_w85, c0_n22_w86, c0_n22_w87, c0_n22_w88, c0_n22_w89, c0_n22_w90, c0_n22_w91, c0_n22_w92, c0_n22_w93, c0_n22_w94, c0_n22_w95, c0_n22_w96, c0_n22_w97, c0_n22_w98, c0_n22_w99, c0_n22_w100, c0_n22_w101, c0_n22_w102, c0_n22_w103, c0_n22_w104, c0_n22_w105, c0_n22_w106, c0_n22_w107, c0_n22_w108, c0_n22_w109, c0_n22_w110, c0_n22_w111, c0_n22_w112, c0_n22_w113, c0_n22_w114, c0_n22_w115, c0_n22_w116, c0_n22_w117, c0_n22_w118, c0_n22_w119, c0_n22_w120, c0_n22_w121, c0_n22_w122, c0_n22_w123, c0_n22_w124, c0_n22_w125, c0_n22_w126, c0_n22_w127, c0_n22_w128, c0_n22_w129, c0_n22_w130, c0_n22_w131, c0_n22_w132, c0_n22_w133, c0_n22_w134, c0_n22_w135, c0_n22_w136, c0_n22_w137, c0_n22_w138, c0_n22_w139, c0_n22_w140, c0_n22_w141, c0_n22_w142, c0_n22_w143, c0_n22_w144, c0_n22_w145, c0_n22_w146, c0_n22_w147, c0_n22_w148, c0_n22_w149, c0_n22_w150, c0_n22_w151, c0_n22_w152, c0_n22_w153, c0_n22_w154, c0_n22_w155, c0_n22_w156, c0_n22_w157, c0_n22_w158, c0_n22_w159, c0_n22_w160, c0_n22_w161, c0_n22_w162, c0_n22_w163, c0_n22_w164, c0_n22_w165, c0_n22_w166, c0_n22_w167, c0_n22_w168, c0_n22_w169, c0_n22_w170, c0_n22_w171, c0_n22_w172, c0_n22_w173, c0_n22_w174, c0_n22_w175, c0_n22_w176, c0_n22_w177, c0_n22_w178, c0_n22_w179, c0_n22_w180, c0_n22_w181, c0_n22_w182, c0_n22_w183, c0_n22_w184, c0_n22_w185, c0_n22_w186, c0_n22_w187, c0_n22_w188, c0_n22_w189, c0_n22_w190, c0_n22_w191, c0_n22_w192, c0_n22_w193, c0_n22_w194, c0_n22_w195, c0_n22_w196, c0_n22_w197, c0_n22_w198, c0_n22_w199, c0_n22_w200, c0_n23_w1, c0_n23_w2, c0_n23_w3, c0_n23_w4, c0_n23_w5, c0_n23_w6, c0_n23_w7, c0_n23_w8, c0_n23_w9, c0_n23_w10, c0_n23_w11, c0_n23_w12, c0_n23_w13, c0_n23_w14, c0_n23_w15, c0_n23_w16, c0_n23_w17, c0_n23_w18, c0_n23_w19, c0_n23_w20, c0_n23_w21, c0_n23_w22, c0_n23_w23, c0_n23_w24, c0_n23_w25, c0_n23_w26, c0_n23_w27, c0_n23_w28, c0_n23_w29, c0_n23_w30, c0_n23_w31, c0_n23_w32, c0_n23_w33, c0_n23_w34, c0_n23_w35, c0_n23_w36, c0_n23_w37, c0_n23_w38, c0_n23_w39, c0_n23_w40, c0_n23_w41, c0_n23_w42, c0_n23_w43, c0_n23_w44, c0_n23_w45, c0_n23_w46, c0_n23_w47, c0_n23_w48, c0_n23_w49, c0_n23_w50, c0_n23_w51, c0_n23_w52, c0_n23_w53, c0_n23_w54, c0_n23_w55, c0_n23_w56, c0_n23_w57, c0_n23_w58, c0_n23_w59, c0_n23_w60, c0_n23_w61, c0_n23_w62, c0_n23_w63, c0_n23_w64, c0_n23_w65, c0_n23_w66, c0_n23_w67, c0_n23_w68, c0_n23_w69, c0_n23_w70, c0_n23_w71, c0_n23_w72, c0_n23_w73, c0_n23_w74, c0_n23_w75, c0_n23_w76, c0_n23_w77, c0_n23_w78, c0_n23_w79, c0_n23_w80, c0_n23_w81, c0_n23_w82, c0_n23_w83, c0_n23_w84, c0_n23_w85, c0_n23_w86, c0_n23_w87, c0_n23_w88, c0_n23_w89, c0_n23_w90, c0_n23_w91, c0_n23_w92, c0_n23_w93, c0_n23_w94, c0_n23_w95, c0_n23_w96, c0_n23_w97, c0_n23_w98, c0_n23_w99, c0_n23_w100, c0_n23_w101, c0_n23_w102, c0_n23_w103, c0_n23_w104, c0_n23_w105, c0_n23_w106, c0_n23_w107, c0_n23_w108, c0_n23_w109, c0_n23_w110, c0_n23_w111, c0_n23_w112, c0_n23_w113, c0_n23_w114, c0_n23_w115, c0_n23_w116, c0_n23_w117, c0_n23_w118, c0_n23_w119, c0_n23_w120, c0_n23_w121, c0_n23_w122, c0_n23_w123, c0_n23_w124, c0_n23_w125, c0_n23_w126, c0_n23_w127, c0_n23_w128, c0_n23_w129, c0_n23_w130, c0_n23_w131, c0_n23_w132, c0_n23_w133, c0_n23_w134, c0_n23_w135, c0_n23_w136, c0_n23_w137, c0_n23_w138, c0_n23_w139, c0_n23_w140, c0_n23_w141, c0_n23_w142, c0_n23_w143, c0_n23_w144, c0_n23_w145, c0_n23_w146, c0_n23_w147, c0_n23_w148, c0_n23_w149, c0_n23_w150, c0_n23_w151, c0_n23_w152, c0_n23_w153, c0_n23_w154, c0_n23_w155, c0_n23_w156, c0_n23_w157, c0_n23_w158, c0_n23_w159, c0_n23_w160, c0_n23_w161, c0_n23_w162, c0_n23_w163, c0_n23_w164, c0_n23_w165, c0_n23_w166, c0_n23_w167, c0_n23_w168, c0_n23_w169, c0_n23_w170, c0_n23_w171, c0_n23_w172, c0_n23_w173, c0_n23_w174, c0_n23_w175, c0_n23_w176, c0_n23_w177, c0_n23_w178, c0_n23_w179, c0_n23_w180, c0_n23_w181, c0_n23_w182, c0_n23_w183, c0_n23_w184, c0_n23_w185, c0_n23_w186, c0_n23_w187, c0_n23_w188, c0_n23_w189, c0_n23_w190, c0_n23_w191, c0_n23_w192, c0_n23_w193, c0_n23_w194, c0_n23_w195, c0_n23_w196, c0_n23_w197, c0_n23_w198, c0_n23_w199, c0_n23_w200, c0_n24_w1, c0_n24_w2, c0_n24_w3, c0_n24_w4, c0_n24_w5, c0_n24_w6, c0_n24_w7, c0_n24_w8, c0_n24_w9, c0_n24_w10, c0_n24_w11, c0_n24_w12, c0_n24_w13, c0_n24_w14, c0_n24_w15, c0_n24_w16, c0_n24_w17, c0_n24_w18, c0_n24_w19, c0_n24_w20, c0_n24_w21, c0_n24_w22, c0_n24_w23, c0_n24_w24, c0_n24_w25, c0_n24_w26, c0_n24_w27, c0_n24_w28, c0_n24_w29, c0_n24_w30, c0_n24_w31, c0_n24_w32, c0_n24_w33, c0_n24_w34, c0_n24_w35, c0_n24_w36, c0_n24_w37, c0_n24_w38, c0_n24_w39, c0_n24_w40, c0_n24_w41, c0_n24_w42, c0_n24_w43, c0_n24_w44, c0_n24_w45, c0_n24_w46, c0_n24_w47, c0_n24_w48, c0_n24_w49, c0_n24_w50, c0_n24_w51, c0_n24_w52, c0_n24_w53, c0_n24_w54, c0_n24_w55, c0_n24_w56, c0_n24_w57, c0_n24_w58, c0_n24_w59, c0_n24_w60, c0_n24_w61, c0_n24_w62, c0_n24_w63, c0_n24_w64, c0_n24_w65, c0_n24_w66, c0_n24_w67, c0_n24_w68, c0_n24_w69, c0_n24_w70, c0_n24_w71, c0_n24_w72, c0_n24_w73, c0_n24_w74, c0_n24_w75, c0_n24_w76, c0_n24_w77, c0_n24_w78, c0_n24_w79, c0_n24_w80, c0_n24_w81, c0_n24_w82, c0_n24_w83, c0_n24_w84, c0_n24_w85, c0_n24_w86, c0_n24_w87, c0_n24_w88, c0_n24_w89, c0_n24_w90, c0_n24_w91, c0_n24_w92, c0_n24_w93, c0_n24_w94, c0_n24_w95, c0_n24_w96, c0_n24_w97, c0_n24_w98, c0_n24_w99, c0_n24_w100, c0_n24_w101, c0_n24_w102, c0_n24_w103, c0_n24_w104, c0_n24_w105, c0_n24_w106, c0_n24_w107, c0_n24_w108, c0_n24_w109, c0_n24_w110, c0_n24_w111, c0_n24_w112, c0_n24_w113, c0_n24_w114, c0_n24_w115, c0_n24_w116, c0_n24_w117, c0_n24_w118, c0_n24_w119, c0_n24_w120, c0_n24_w121, c0_n24_w122, c0_n24_w123, c0_n24_w124, c0_n24_w125, c0_n24_w126, c0_n24_w127, c0_n24_w128, c0_n24_w129, c0_n24_w130, c0_n24_w131, c0_n24_w132, c0_n24_w133, c0_n24_w134, c0_n24_w135, c0_n24_w136, c0_n24_w137, c0_n24_w138, c0_n24_w139, c0_n24_w140, c0_n24_w141, c0_n24_w142, c0_n24_w143, c0_n24_w144, c0_n24_w145, c0_n24_w146, c0_n24_w147, c0_n24_w148, c0_n24_w149, c0_n24_w150, c0_n24_w151, c0_n24_w152, c0_n24_w153, c0_n24_w154, c0_n24_w155, c0_n24_w156, c0_n24_w157, c0_n24_w158, c0_n24_w159, c0_n24_w160, c0_n24_w161, c0_n24_w162, c0_n24_w163, c0_n24_w164, c0_n24_w165, c0_n24_w166, c0_n24_w167, c0_n24_w168, c0_n24_w169, c0_n24_w170, c0_n24_w171, c0_n24_w172, c0_n24_w173, c0_n24_w174, c0_n24_w175, c0_n24_w176, c0_n24_w177, c0_n24_w178, c0_n24_w179, c0_n24_w180, c0_n24_w181, c0_n24_w182, c0_n24_w183, c0_n24_w184, c0_n24_w185, c0_n24_w186, c0_n24_w187, c0_n24_w188, c0_n24_w189, c0_n24_w190, c0_n24_w191, c0_n24_w192, c0_n24_w193, c0_n24_w194, c0_n24_w195, c0_n24_w196, c0_n24_w197, c0_n24_w198, c0_n24_w199, c0_n24_w200, c0_n25_w1, c0_n25_w2, c0_n25_w3, c0_n25_w4, c0_n25_w5, c0_n25_w6, c0_n25_w7, c0_n25_w8, c0_n25_w9, c0_n25_w10, c0_n25_w11, c0_n25_w12, c0_n25_w13, c0_n25_w14, c0_n25_w15, c0_n25_w16, c0_n25_w17, c0_n25_w18, c0_n25_w19, c0_n25_w20, c0_n25_w21, c0_n25_w22, c0_n25_w23, c0_n25_w24, c0_n25_w25, c0_n25_w26, c0_n25_w27, c0_n25_w28, c0_n25_w29, c0_n25_w30, c0_n25_w31, c0_n25_w32, c0_n25_w33, c0_n25_w34, c0_n25_w35, c0_n25_w36, c0_n25_w37, c0_n25_w38, c0_n25_w39, c0_n25_w40, c0_n25_w41, c0_n25_w42, c0_n25_w43, c0_n25_w44, c0_n25_w45, c0_n25_w46, c0_n25_w47, c0_n25_w48, c0_n25_w49, c0_n25_w50, c0_n25_w51, c0_n25_w52, c0_n25_w53, c0_n25_w54, c0_n25_w55, c0_n25_w56, c0_n25_w57, c0_n25_w58, c0_n25_w59, c0_n25_w60, c0_n25_w61, c0_n25_w62, c0_n25_w63, c0_n25_w64, c0_n25_w65, c0_n25_w66, c0_n25_w67, c0_n25_w68, c0_n25_w69, c0_n25_w70, c0_n25_w71, c0_n25_w72, c0_n25_w73, c0_n25_w74, c0_n25_w75, c0_n25_w76, c0_n25_w77, c0_n25_w78, c0_n25_w79, c0_n25_w80, c0_n25_w81, c0_n25_w82, c0_n25_w83, c0_n25_w84, c0_n25_w85, c0_n25_w86, c0_n25_w87, c0_n25_w88, c0_n25_w89, c0_n25_w90, c0_n25_w91, c0_n25_w92, c0_n25_w93, c0_n25_w94, c0_n25_w95, c0_n25_w96, c0_n25_w97, c0_n25_w98, c0_n25_w99, c0_n25_w100, c0_n25_w101, c0_n25_w102, c0_n25_w103, c0_n25_w104, c0_n25_w105, c0_n25_w106, c0_n25_w107, c0_n25_w108, c0_n25_w109, c0_n25_w110, c0_n25_w111, c0_n25_w112, c0_n25_w113, c0_n25_w114, c0_n25_w115, c0_n25_w116, c0_n25_w117, c0_n25_w118, c0_n25_w119, c0_n25_w120, c0_n25_w121, c0_n25_w122, c0_n25_w123, c0_n25_w124, c0_n25_w125, c0_n25_w126, c0_n25_w127, c0_n25_w128, c0_n25_w129, c0_n25_w130, c0_n25_w131, c0_n25_w132, c0_n25_w133, c0_n25_w134, c0_n25_w135, c0_n25_w136, c0_n25_w137, c0_n25_w138, c0_n25_w139, c0_n25_w140, c0_n25_w141, c0_n25_w142, c0_n25_w143, c0_n25_w144, c0_n25_w145, c0_n25_w146, c0_n25_w147, c0_n25_w148, c0_n25_w149, c0_n25_w150, c0_n25_w151, c0_n25_w152, c0_n25_w153, c0_n25_w154, c0_n25_w155, c0_n25_w156, c0_n25_w157, c0_n25_w158, c0_n25_w159, c0_n25_w160, c0_n25_w161, c0_n25_w162, c0_n25_w163, c0_n25_w164, c0_n25_w165, c0_n25_w166, c0_n25_w167, c0_n25_w168, c0_n25_w169, c0_n25_w170, c0_n25_w171, c0_n25_w172, c0_n25_w173, c0_n25_w174, c0_n25_w175, c0_n25_w176, c0_n25_w177, c0_n25_w178, c0_n25_w179, c0_n25_w180, c0_n25_w181, c0_n25_w182, c0_n25_w183, c0_n25_w184, c0_n25_w185, c0_n25_w186, c0_n25_w187, c0_n25_w188, c0_n25_w189, c0_n25_w190, c0_n25_w191, c0_n25_w192, c0_n25_w193, c0_n25_w194, c0_n25_w195, c0_n25_w196, c0_n25_w197, c0_n25_w198, c0_n25_w199, c0_n25_w200, c0_n26_w1, c0_n26_w2, c0_n26_w3, c0_n26_w4, c0_n26_w5, c0_n26_w6, c0_n26_w7, c0_n26_w8, c0_n26_w9, c0_n26_w10, c0_n26_w11, c0_n26_w12, c0_n26_w13, c0_n26_w14, c0_n26_w15, c0_n26_w16, c0_n26_w17, c0_n26_w18, c0_n26_w19, c0_n26_w20, c0_n26_w21, c0_n26_w22, c0_n26_w23, c0_n26_w24, c0_n26_w25, c0_n26_w26, c0_n26_w27, c0_n26_w28, c0_n26_w29, c0_n26_w30, c0_n26_w31, c0_n26_w32, c0_n26_w33, c0_n26_w34, c0_n26_w35, c0_n26_w36, c0_n26_w37, c0_n26_w38, c0_n26_w39, c0_n26_w40, c0_n26_w41, c0_n26_w42, c0_n26_w43, c0_n26_w44, c0_n26_w45, c0_n26_w46, c0_n26_w47, c0_n26_w48, c0_n26_w49, c0_n26_w50, c0_n26_w51, c0_n26_w52, c0_n26_w53, c0_n26_w54, c0_n26_w55, c0_n26_w56, c0_n26_w57, c0_n26_w58, c0_n26_w59, c0_n26_w60, c0_n26_w61, c0_n26_w62, c0_n26_w63, c0_n26_w64, c0_n26_w65, c0_n26_w66, c0_n26_w67, c0_n26_w68, c0_n26_w69, c0_n26_w70, c0_n26_w71, c0_n26_w72, c0_n26_w73, c0_n26_w74, c0_n26_w75, c0_n26_w76, c0_n26_w77, c0_n26_w78, c0_n26_w79, c0_n26_w80, c0_n26_w81, c0_n26_w82, c0_n26_w83, c0_n26_w84, c0_n26_w85, c0_n26_w86, c0_n26_w87, c0_n26_w88, c0_n26_w89, c0_n26_w90, c0_n26_w91, c0_n26_w92, c0_n26_w93, c0_n26_w94, c0_n26_w95, c0_n26_w96, c0_n26_w97, c0_n26_w98, c0_n26_w99, c0_n26_w100, c0_n26_w101, c0_n26_w102, c0_n26_w103, c0_n26_w104, c0_n26_w105, c0_n26_w106, c0_n26_w107, c0_n26_w108, c0_n26_w109, c0_n26_w110, c0_n26_w111, c0_n26_w112, c0_n26_w113, c0_n26_w114, c0_n26_w115, c0_n26_w116, c0_n26_w117, c0_n26_w118, c0_n26_w119, c0_n26_w120, c0_n26_w121, c0_n26_w122, c0_n26_w123, c0_n26_w124, c0_n26_w125, c0_n26_w126, c0_n26_w127, c0_n26_w128, c0_n26_w129, c0_n26_w130, c0_n26_w131, c0_n26_w132, c0_n26_w133, c0_n26_w134, c0_n26_w135, c0_n26_w136, c0_n26_w137, c0_n26_w138, c0_n26_w139, c0_n26_w140, c0_n26_w141, c0_n26_w142, c0_n26_w143, c0_n26_w144, c0_n26_w145, c0_n26_w146, c0_n26_w147, c0_n26_w148, c0_n26_w149, c0_n26_w150, c0_n26_w151, c0_n26_w152, c0_n26_w153, c0_n26_w154, c0_n26_w155, c0_n26_w156, c0_n26_w157, c0_n26_w158, c0_n26_w159, c0_n26_w160, c0_n26_w161, c0_n26_w162, c0_n26_w163, c0_n26_w164, c0_n26_w165, c0_n26_w166, c0_n26_w167, c0_n26_w168, c0_n26_w169, c0_n26_w170, c0_n26_w171, c0_n26_w172, c0_n26_w173, c0_n26_w174, c0_n26_w175, c0_n26_w176, c0_n26_w177, c0_n26_w178, c0_n26_w179, c0_n26_w180, c0_n26_w181, c0_n26_w182, c0_n26_w183, c0_n26_w184, c0_n26_w185, c0_n26_w186, c0_n26_w187, c0_n26_w188, c0_n26_w189, c0_n26_w190, c0_n26_w191, c0_n26_w192, c0_n26_w193, c0_n26_w194, c0_n26_w195, c0_n26_w196, c0_n26_w197, c0_n26_w198, c0_n26_w199, c0_n26_w200, c0_n27_w1, c0_n27_w2, c0_n27_w3, c0_n27_w4, c0_n27_w5, c0_n27_w6, c0_n27_w7, c0_n27_w8, c0_n27_w9, c0_n27_w10, c0_n27_w11, c0_n27_w12, c0_n27_w13, c0_n27_w14, c0_n27_w15, c0_n27_w16, c0_n27_w17, c0_n27_w18, c0_n27_w19, c0_n27_w20, c0_n27_w21, c0_n27_w22, c0_n27_w23, c0_n27_w24, c0_n27_w25, c0_n27_w26, c0_n27_w27, c0_n27_w28, c0_n27_w29, c0_n27_w30, c0_n27_w31, c0_n27_w32, c0_n27_w33, c0_n27_w34, c0_n27_w35, c0_n27_w36, c0_n27_w37, c0_n27_w38, c0_n27_w39, c0_n27_w40, c0_n27_w41, c0_n27_w42, c0_n27_w43, c0_n27_w44, c0_n27_w45, c0_n27_w46, c0_n27_w47, c0_n27_w48, c0_n27_w49, c0_n27_w50, c0_n27_w51, c0_n27_w52, c0_n27_w53, c0_n27_w54, c0_n27_w55, c0_n27_w56, c0_n27_w57, c0_n27_w58, c0_n27_w59, c0_n27_w60, c0_n27_w61, c0_n27_w62, c0_n27_w63, c0_n27_w64, c0_n27_w65, c0_n27_w66, c0_n27_w67, c0_n27_w68, c0_n27_w69, c0_n27_w70, c0_n27_w71, c0_n27_w72, c0_n27_w73, c0_n27_w74, c0_n27_w75, c0_n27_w76, c0_n27_w77, c0_n27_w78, c0_n27_w79, c0_n27_w80, c0_n27_w81, c0_n27_w82, c0_n27_w83, c0_n27_w84, c0_n27_w85, c0_n27_w86, c0_n27_w87, c0_n27_w88, c0_n27_w89, c0_n27_w90, c0_n27_w91, c0_n27_w92, c0_n27_w93, c0_n27_w94, c0_n27_w95, c0_n27_w96, c0_n27_w97, c0_n27_w98, c0_n27_w99, c0_n27_w100, c0_n27_w101, c0_n27_w102, c0_n27_w103, c0_n27_w104, c0_n27_w105, c0_n27_w106, c0_n27_w107, c0_n27_w108, c0_n27_w109, c0_n27_w110, c0_n27_w111, c0_n27_w112, c0_n27_w113, c0_n27_w114, c0_n27_w115, c0_n27_w116, c0_n27_w117, c0_n27_w118, c0_n27_w119, c0_n27_w120, c0_n27_w121, c0_n27_w122, c0_n27_w123, c0_n27_w124, c0_n27_w125, c0_n27_w126, c0_n27_w127, c0_n27_w128, c0_n27_w129, c0_n27_w130, c0_n27_w131, c0_n27_w132, c0_n27_w133, c0_n27_w134, c0_n27_w135, c0_n27_w136, c0_n27_w137, c0_n27_w138, c0_n27_w139, c0_n27_w140, c0_n27_w141, c0_n27_w142, c0_n27_w143, c0_n27_w144, c0_n27_w145, c0_n27_w146, c0_n27_w147, c0_n27_w148, c0_n27_w149, c0_n27_w150, c0_n27_w151, c0_n27_w152, c0_n27_w153, c0_n27_w154, c0_n27_w155, c0_n27_w156, c0_n27_w157, c0_n27_w158, c0_n27_w159, c0_n27_w160, c0_n27_w161, c0_n27_w162, c0_n27_w163, c0_n27_w164, c0_n27_w165, c0_n27_w166, c0_n27_w167, c0_n27_w168, c0_n27_w169, c0_n27_w170, c0_n27_w171, c0_n27_w172, c0_n27_w173, c0_n27_w174, c0_n27_w175, c0_n27_w176, c0_n27_w177, c0_n27_w178, c0_n27_w179, c0_n27_w180, c0_n27_w181, c0_n27_w182, c0_n27_w183, c0_n27_w184, c0_n27_w185, c0_n27_w186, c0_n27_w187, c0_n27_w188, c0_n27_w189, c0_n27_w190, c0_n27_w191, c0_n27_w192, c0_n27_w193, c0_n27_w194, c0_n27_w195, c0_n27_w196, c0_n27_w197, c0_n27_w198, c0_n27_w199, c0_n27_w200, c0_n28_w1, c0_n28_w2, c0_n28_w3, c0_n28_w4, c0_n28_w5, c0_n28_w6, c0_n28_w7, c0_n28_w8, c0_n28_w9, c0_n28_w10, c0_n28_w11, c0_n28_w12, c0_n28_w13, c0_n28_w14, c0_n28_w15, c0_n28_w16, c0_n28_w17, c0_n28_w18, c0_n28_w19, c0_n28_w20, c0_n28_w21, c0_n28_w22, c0_n28_w23, c0_n28_w24, c0_n28_w25, c0_n28_w26, c0_n28_w27, c0_n28_w28, c0_n28_w29, c0_n28_w30, c0_n28_w31, c0_n28_w32, c0_n28_w33, c0_n28_w34, c0_n28_w35, c0_n28_w36, c0_n28_w37, c0_n28_w38, c0_n28_w39, c0_n28_w40, c0_n28_w41, c0_n28_w42, c0_n28_w43, c0_n28_w44, c0_n28_w45, c0_n28_w46, c0_n28_w47, c0_n28_w48, c0_n28_w49, c0_n28_w50, c0_n28_w51, c0_n28_w52, c0_n28_w53, c0_n28_w54, c0_n28_w55, c0_n28_w56, c0_n28_w57, c0_n28_w58, c0_n28_w59, c0_n28_w60, c0_n28_w61, c0_n28_w62, c0_n28_w63, c0_n28_w64, c0_n28_w65, c0_n28_w66, c0_n28_w67, c0_n28_w68, c0_n28_w69, c0_n28_w70, c0_n28_w71, c0_n28_w72, c0_n28_w73, c0_n28_w74, c0_n28_w75, c0_n28_w76, c0_n28_w77, c0_n28_w78, c0_n28_w79, c0_n28_w80, c0_n28_w81, c0_n28_w82, c0_n28_w83, c0_n28_w84, c0_n28_w85, c0_n28_w86, c0_n28_w87, c0_n28_w88, c0_n28_w89, c0_n28_w90, c0_n28_w91, c0_n28_w92, c0_n28_w93, c0_n28_w94, c0_n28_w95, c0_n28_w96, c0_n28_w97, c0_n28_w98, c0_n28_w99, c0_n28_w100, c0_n28_w101, c0_n28_w102, c0_n28_w103, c0_n28_w104, c0_n28_w105, c0_n28_w106, c0_n28_w107, c0_n28_w108, c0_n28_w109, c0_n28_w110, c0_n28_w111, c0_n28_w112, c0_n28_w113, c0_n28_w114, c0_n28_w115, c0_n28_w116, c0_n28_w117, c0_n28_w118, c0_n28_w119, c0_n28_w120, c0_n28_w121, c0_n28_w122, c0_n28_w123, c0_n28_w124, c0_n28_w125, c0_n28_w126, c0_n28_w127, c0_n28_w128, c0_n28_w129, c0_n28_w130, c0_n28_w131, c0_n28_w132, c0_n28_w133, c0_n28_w134, c0_n28_w135, c0_n28_w136, c0_n28_w137, c0_n28_w138, c0_n28_w139, c0_n28_w140, c0_n28_w141, c0_n28_w142, c0_n28_w143, c0_n28_w144, c0_n28_w145, c0_n28_w146, c0_n28_w147, c0_n28_w148, c0_n28_w149, c0_n28_w150, c0_n28_w151, c0_n28_w152, c0_n28_w153, c0_n28_w154, c0_n28_w155, c0_n28_w156, c0_n28_w157, c0_n28_w158, c0_n28_w159, c0_n28_w160, c0_n28_w161, c0_n28_w162, c0_n28_w163, c0_n28_w164, c0_n28_w165, c0_n28_w166, c0_n28_w167, c0_n28_w168, c0_n28_w169, c0_n28_w170, c0_n28_w171, c0_n28_w172, c0_n28_w173, c0_n28_w174, c0_n28_w175, c0_n28_w176, c0_n28_w177, c0_n28_w178, c0_n28_w179, c0_n28_w180, c0_n28_w181, c0_n28_w182, c0_n28_w183, c0_n28_w184, c0_n28_w185, c0_n28_w186, c0_n28_w187, c0_n28_w188, c0_n28_w189, c0_n28_w190, c0_n28_w191, c0_n28_w192, c0_n28_w193, c0_n28_w194, c0_n28_w195, c0_n28_w196, c0_n28_w197, c0_n28_w198, c0_n28_w199, c0_n28_w200, c0_n29_w1, c0_n29_w2, c0_n29_w3, c0_n29_w4, c0_n29_w5, c0_n29_w6, c0_n29_w7, c0_n29_w8, c0_n29_w9, c0_n29_w10, c0_n29_w11, c0_n29_w12, c0_n29_w13, c0_n29_w14, c0_n29_w15, c0_n29_w16, c0_n29_w17, c0_n29_w18, c0_n29_w19, c0_n29_w20, c0_n29_w21, c0_n29_w22, c0_n29_w23, c0_n29_w24, c0_n29_w25, c0_n29_w26, c0_n29_w27, c0_n29_w28, c0_n29_w29, c0_n29_w30, c0_n29_w31, c0_n29_w32, c0_n29_w33, c0_n29_w34, c0_n29_w35, c0_n29_w36, c0_n29_w37, c0_n29_w38, c0_n29_w39, c0_n29_w40, c0_n29_w41, c0_n29_w42, c0_n29_w43, c0_n29_w44, c0_n29_w45, c0_n29_w46, c0_n29_w47, c0_n29_w48, c0_n29_w49, c0_n29_w50, c0_n29_w51, c0_n29_w52, c0_n29_w53, c0_n29_w54, c0_n29_w55, c0_n29_w56, c0_n29_w57, c0_n29_w58, c0_n29_w59, c0_n29_w60, c0_n29_w61, c0_n29_w62, c0_n29_w63, c0_n29_w64, c0_n29_w65, c0_n29_w66, c0_n29_w67, c0_n29_w68, c0_n29_w69, c0_n29_w70, c0_n29_w71, c0_n29_w72, c0_n29_w73, c0_n29_w74, c0_n29_w75, c0_n29_w76, c0_n29_w77, c0_n29_w78, c0_n29_w79, c0_n29_w80, c0_n29_w81, c0_n29_w82, c0_n29_w83, c0_n29_w84, c0_n29_w85, c0_n29_w86, c0_n29_w87, c0_n29_w88, c0_n29_w89, c0_n29_w90, c0_n29_w91, c0_n29_w92, c0_n29_w93, c0_n29_w94, c0_n29_w95, c0_n29_w96, c0_n29_w97, c0_n29_w98, c0_n29_w99, c0_n29_w100, c0_n29_w101, c0_n29_w102, c0_n29_w103, c0_n29_w104, c0_n29_w105, c0_n29_w106, c0_n29_w107, c0_n29_w108, c0_n29_w109, c0_n29_w110, c0_n29_w111, c0_n29_w112, c0_n29_w113, c0_n29_w114, c0_n29_w115, c0_n29_w116, c0_n29_w117, c0_n29_w118, c0_n29_w119, c0_n29_w120, c0_n29_w121, c0_n29_w122, c0_n29_w123, c0_n29_w124, c0_n29_w125, c0_n29_w126, c0_n29_w127, c0_n29_w128, c0_n29_w129, c0_n29_w130, c0_n29_w131, c0_n29_w132, c0_n29_w133, c0_n29_w134, c0_n29_w135, c0_n29_w136, c0_n29_w137, c0_n29_w138, c0_n29_w139, c0_n29_w140, c0_n29_w141, c0_n29_w142, c0_n29_w143, c0_n29_w144, c0_n29_w145, c0_n29_w146, c0_n29_w147, c0_n29_w148, c0_n29_w149, c0_n29_w150, c0_n29_w151, c0_n29_w152, c0_n29_w153, c0_n29_w154, c0_n29_w155, c0_n29_w156, c0_n29_w157, c0_n29_w158, c0_n29_w159, c0_n29_w160, c0_n29_w161, c0_n29_w162, c0_n29_w163, c0_n29_w164, c0_n29_w165, c0_n29_w166, c0_n29_w167, c0_n29_w168, c0_n29_w169, c0_n29_w170, c0_n29_w171, c0_n29_w172, c0_n29_w173, c0_n29_w174, c0_n29_w175, c0_n29_w176, c0_n29_w177, c0_n29_w178, c0_n29_w179, c0_n29_w180, c0_n29_w181, c0_n29_w182, c0_n29_w183, c0_n29_w184, c0_n29_w185, c0_n29_w186, c0_n29_w187, c0_n29_w188, c0_n29_w189, c0_n29_w190, c0_n29_w191, c0_n29_w192, c0_n29_w193, c0_n29_w194, c0_n29_w195, c0_n29_w196, c0_n29_w197, c0_n29_w198, c0_n29_w199, c0_n29_w200, c0_n30_w1, c0_n30_w2, c0_n30_w3, c0_n30_w4, c0_n30_w5, c0_n30_w6, c0_n30_w7, c0_n30_w8, c0_n30_w9, c0_n30_w10, c0_n30_w11, c0_n30_w12, c0_n30_w13, c0_n30_w14, c0_n30_w15, c0_n30_w16, c0_n30_w17, c0_n30_w18, c0_n30_w19, c0_n30_w20, c0_n30_w21, c0_n30_w22, c0_n30_w23, c0_n30_w24, c0_n30_w25, c0_n30_w26, c0_n30_w27, c0_n30_w28, c0_n30_w29, c0_n30_w30, c0_n30_w31, c0_n30_w32, c0_n30_w33, c0_n30_w34, c0_n30_w35, c0_n30_w36, c0_n30_w37, c0_n30_w38, c0_n30_w39, c0_n30_w40, c0_n30_w41, c0_n30_w42, c0_n30_w43, c0_n30_w44, c0_n30_w45, c0_n30_w46, c0_n30_w47, c0_n30_w48, c0_n30_w49, c0_n30_w50, c0_n30_w51, c0_n30_w52, c0_n30_w53, c0_n30_w54, c0_n30_w55, c0_n30_w56, c0_n30_w57, c0_n30_w58, c0_n30_w59, c0_n30_w60, c0_n30_w61, c0_n30_w62, c0_n30_w63, c0_n30_w64, c0_n30_w65, c0_n30_w66, c0_n30_w67, c0_n30_w68, c0_n30_w69, c0_n30_w70, c0_n30_w71, c0_n30_w72, c0_n30_w73, c0_n30_w74, c0_n30_w75, c0_n30_w76, c0_n30_w77, c0_n30_w78, c0_n30_w79, c0_n30_w80, c0_n30_w81, c0_n30_w82, c0_n30_w83, c0_n30_w84, c0_n30_w85, c0_n30_w86, c0_n30_w87, c0_n30_w88, c0_n30_w89, c0_n30_w90, c0_n30_w91, c0_n30_w92, c0_n30_w93, c0_n30_w94, c0_n30_w95, c0_n30_w96, c0_n30_w97, c0_n30_w98, c0_n30_w99, c0_n30_w100, c0_n30_w101, c0_n30_w102, c0_n30_w103, c0_n30_w104, c0_n30_w105, c0_n30_w106, c0_n30_w107, c0_n30_w108, c0_n30_w109, c0_n30_w110, c0_n30_w111, c0_n30_w112, c0_n30_w113, c0_n30_w114, c0_n30_w115, c0_n30_w116, c0_n30_w117, c0_n30_w118, c0_n30_w119, c0_n30_w120, c0_n30_w121, c0_n30_w122, c0_n30_w123, c0_n30_w124, c0_n30_w125, c0_n30_w126, c0_n30_w127, c0_n30_w128, c0_n30_w129, c0_n30_w130, c0_n30_w131, c0_n30_w132, c0_n30_w133, c0_n30_w134, c0_n30_w135, c0_n30_w136, c0_n30_w137, c0_n30_w138, c0_n30_w139, c0_n30_w140, c0_n30_w141, c0_n30_w142, c0_n30_w143, c0_n30_w144, c0_n30_w145, c0_n30_w146, c0_n30_w147, c0_n30_w148, c0_n30_w149, c0_n30_w150, c0_n30_w151, c0_n30_w152, c0_n30_w153, c0_n30_w154, c0_n30_w155, c0_n30_w156, c0_n30_w157, c0_n30_w158, c0_n30_w159, c0_n30_w160, c0_n30_w161, c0_n30_w162, c0_n30_w163, c0_n30_w164, c0_n30_w165, c0_n30_w166, c0_n30_w167, c0_n30_w168, c0_n30_w169, c0_n30_w170, c0_n30_w171, c0_n30_w172, c0_n30_w173, c0_n30_w174, c0_n30_w175, c0_n30_w176, c0_n30_w177, c0_n30_w178, c0_n30_w179, c0_n30_w180, c0_n30_w181, c0_n30_w182, c0_n30_w183, c0_n30_w184, c0_n30_w185, c0_n30_w186, c0_n30_w187, c0_n30_w188, c0_n30_w189, c0_n30_w190, c0_n30_w191, c0_n30_w192, c0_n30_w193, c0_n30_w194, c0_n30_w195, c0_n30_w196, c0_n30_w197, c0_n30_w198, c0_n30_w199, c0_n30_w200, c0_n31_w1, c0_n31_w2, c0_n31_w3, c0_n31_w4, c0_n31_w5, c0_n31_w6, c0_n31_w7, c0_n31_w8, c0_n31_w9, c0_n31_w10, c0_n31_w11, c0_n31_w12, c0_n31_w13, c0_n31_w14, c0_n31_w15, c0_n31_w16, c0_n31_w17, c0_n31_w18, c0_n31_w19, c0_n31_w20, c0_n31_w21, c0_n31_w22, c0_n31_w23, c0_n31_w24, c0_n31_w25, c0_n31_w26, c0_n31_w27, c0_n31_w28, c0_n31_w29, c0_n31_w30, c0_n31_w31, c0_n31_w32, c0_n31_w33, c0_n31_w34, c0_n31_w35, c0_n31_w36, c0_n31_w37, c0_n31_w38, c0_n31_w39, c0_n31_w40, c0_n31_w41, c0_n31_w42, c0_n31_w43, c0_n31_w44, c0_n31_w45, c0_n31_w46, c0_n31_w47, c0_n31_w48, c0_n31_w49, c0_n31_w50, c0_n31_w51, c0_n31_w52, c0_n31_w53, c0_n31_w54, c0_n31_w55, c0_n31_w56, c0_n31_w57, c0_n31_w58, c0_n31_w59, c0_n31_w60, c0_n31_w61, c0_n31_w62, c0_n31_w63, c0_n31_w64, c0_n31_w65, c0_n31_w66, c0_n31_w67, c0_n31_w68, c0_n31_w69, c0_n31_w70, c0_n31_w71, c0_n31_w72, c0_n31_w73, c0_n31_w74, c0_n31_w75, c0_n31_w76, c0_n31_w77, c0_n31_w78, c0_n31_w79, c0_n31_w80, c0_n31_w81, c0_n31_w82, c0_n31_w83, c0_n31_w84, c0_n31_w85, c0_n31_w86, c0_n31_w87, c0_n31_w88, c0_n31_w89, c0_n31_w90, c0_n31_w91, c0_n31_w92, c0_n31_w93, c0_n31_w94, c0_n31_w95, c0_n31_w96, c0_n31_w97, c0_n31_w98, c0_n31_w99, c0_n31_w100, c0_n31_w101, c0_n31_w102, c0_n31_w103, c0_n31_w104, c0_n31_w105, c0_n31_w106, c0_n31_w107, c0_n31_w108, c0_n31_w109, c0_n31_w110, c0_n31_w111, c0_n31_w112, c0_n31_w113, c0_n31_w114, c0_n31_w115, c0_n31_w116, c0_n31_w117, c0_n31_w118, c0_n31_w119, c0_n31_w120, c0_n31_w121, c0_n31_w122, c0_n31_w123, c0_n31_w124, c0_n31_w125, c0_n31_w126, c0_n31_w127, c0_n31_w128, c0_n31_w129, c0_n31_w130, c0_n31_w131, c0_n31_w132, c0_n31_w133, c0_n31_w134, c0_n31_w135, c0_n31_w136, c0_n31_w137, c0_n31_w138, c0_n31_w139, c0_n31_w140, c0_n31_w141, c0_n31_w142, c0_n31_w143, c0_n31_w144, c0_n31_w145, c0_n31_w146, c0_n31_w147, c0_n31_w148, c0_n31_w149, c0_n31_w150, c0_n31_w151, c0_n31_w152, c0_n31_w153, c0_n31_w154, c0_n31_w155, c0_n31_w156, c0_n31_w157, c0_n31_w158, c0_n31_w159, c0_n31_w160, c0_n31_w161, c0_n31_w162, c0_n31_w163, c0_n31_w164, c0_n31_w165, c0_n31_w166, c0_n31_w167, c0_n31_w168, c0_n31_w169, c0_n31_w170, c0_n31_w171, c0_n31_w172, c0_n31_w173, c0_n31_w174, c0_n31_w175, c0_n31_w176, c0_n31_w177, c0_n31_w178, c0_n31_w179, c0_n31_w180, c0_n31_w181, c0_n31_w182, c0_n31_w183, c0_n31_w184, c0_n31_w185, c0_n31_w186, c0_n31_w187, c0_n31_w188, c0_n31_w189, c0_n31_w190, c0_n31_w191, c0_n31_w192, c0_n31_w193, c0_n31_w194, c0_n31_w195, c0_n31_w196, c0_n31_w197, c0_n31_w198, c0_n31_w199, c0_n31_w200, c0_n32_w1, c0_n32_w2, c0_n32_w3, c0_n32_w4, c0_n32_w5, c0_n32_w6, c0_n32_w7, c0_n32_w8, c0_n32_w9, c0_n32_w10, c0_n32_w11, c0_n32_w12, c0_n32_w13, c0_n32_w14, c0_n32_w15, c0_n32_w16, c0_n32_w17, c0_n32_w18, c0_n32_w19, c0_n32_w20, c0_n32_w21, c0_n32_w22, c0_n32_w23, c0_n32_w24, c0_n32_w25, c0_n32_w26, c0_n32_w27, c0_n32_w28, c0_n32_w29, c0_n32_w30, c0_n32_w31, c0_n32_w32, c0_n32_w33, c0_n32_w34, c0_n32_w35, c0_n32_w36, c0_n32_w37, c0_n32_w38, c0_n32_w39, c0_n32_w40, c0_n32_w41, c0_n32_w42, c0_n32_w43, c0_n32_w44, c0_n32_w45, c0_n32_w46, c0_n32_w47, c0_n32_w48, c0_n32_w49, c0_n32_w50, c0_n32_w51, c0_n32_w52, c0_n32_w53, c0_n32_w54, c0_n32_w55, c0_n32_w56, c0_n32_w57, c0_n32_w58, c0_n32_w59, c0_n32_w60, c0_n32_w61, c0_n32_w62, c0_n32_w63, c0_n32_w64, c0_n32_w65, c0_n32_w66, c0_n32_w67, c0_n32_w68, c0_n32_w69, c0_n32_w70, c0_n32_w71, c0_n32_w72, c0_n32_w73, c0_n32_w74, c0_n32_w75, c0_n32_w76, c0_n32_w77, c0_n32_w78, c0_n32_w79, c0_n32_w80, c0_n32_w81, c0_n32_w82, c0_n32_w83, c0_n32_w84, c0_n32_w85, c0_n32_w86, c0_n32_w87, c0_n32_w88, c0_n32_w89, c0_n32_w90, c0_n32_w91, c0_n32_w92, c0_n32_w93, c0_n32_w94, c0_n32_w95, c0_n32_w96, c0_n32_w97, c0_n32_w98, c0_n32_w99, c0_n32_w100, c0_n32_w101, c0_n32_w102, c0_n32_w103, c0_n32_w104, c0_n32_w105, c0_n32_w106, c0_n32_w107, c0_n32_w108, c0_n32_w109, c0_n32_w110, c0_n32_w111, c0_n32_w112, c0_n32_w113, c0_n32_w114, c0_n32_w115, c0_n32_w116, c0_n32_w117, c0_n32_w118, c0_n32_w119, c0_n32_w120, c0_n32_w121, c0_n32_w122, c0_n32_w123, c0_n32_w124, c0_n32_w125, c0_n32_w126, c0_n32_w127, c0_n32_w128, c0_n32_w129, c0_n32_w130, c0_n32_w131, c0_n32_w132, c0_n32_w133, c0_n32_w134, c0_n32_w135, c0_n32_w136, c0_n32_w137, c0_n32_w138, c0_n32_w139, c0_n32_w140, c0_n32_w141, c0_n32_w142, c0_n32_w143, c0_n32_w144, c0_n32_w145, c0_n32_w146, c0_n32_w147, c0_n32_w148, c0_n32_w149, c0_n32_w150, c0_n32_w151, c0_n32_w152, c0_n32_w153, c0_n32_w154, c0_n32_w155, c0_n32_w156, c0_n32_w157, c0_n32_w158, c0_n32_w159, c0_n32_w160, c0_n32_w161, c0_n32_w162, c0_n32_w163, c0_n32_w164, c0_n32_w165, c0_n32_w166, c0_n32_w167, c0_n32_w168, c0_n32_w169, c0_n32_w170, c0_n32_w171, c0_n32_w172, c0_n32_w173, c0_n32_w174, c0_n32_w175, c0_n32_w176, c0_n32_w177, c0_n32_w178, c0_n32_w179, c0_n32_w180, c0_n32_w181, c0_n32_w182, c0_n32_w183, c0_n32_w184, c0_n32_w185, c0_n32_w186, c0_n32_w187, c0_n32_w188, c0_n32_w189, c0_n32_w190, c0_n32_w191, c0_n32_w192, c0_n32_w193, c0_n32_w194, c0_n32_w195, c0_n32_w196, c0_n32_w197, c0_n32_w198, c0_n32_w199, c0_n32_w200, c0_n33_w1, c0_n33_w2, c0_n33_w3, c0_n33_w4, c0_n33_w5, c0_n33_w6, c0_n33_w7, c0_n33_w8, c0_n33_w9, c0_n33_w10, c0_n33_w11, c0_n33_w12, c0_n33_w13, c0_n33_w14, c0_n33_w15, c0_n33_w16, c0_n33_w17, c0_n33_w18, c0_n33_w19, c0_n33_w20, c0_n33_w21, c0_n33_w22, c0_n33_w23, c0_n33_w24, c0_n33_w25, c0_n33_w26, c0_n33_w27, c0_n33_w28, c0_n33_w29, c0_n33_w30, c0_n33_w31, c0_n33_w32, c0_n33_w33, c0_n33_w34, c0_n33_w35, c0_n33_w36, c0_n33_w37, c0_n33_w38, c0_n33_w39, c0_n33_w40, c0_n33_w41, c0_n33_w42, c0_n33_w43, c0_n33_w44, c0_n33_w45, c0_n33_w46, c0_n33_w47, c0_n33_w48, c0_n33_w49, c0_n33_w50, c0_n33_w51, c0_n33_w52, c0_n33_w53, c0_n33_w54, c0_n33_w55, c0_n33_w56, c0_n33_w57, c0_n33_w58, c0_n33_w59, c0_n33_w60, c0_n33_w61, c0_n33_w62, c0_n33_w63, c0_n33_w64, c0_n33_w65, c0_n33_w66, c0_n33_w67, c0_n33_w68, c0_n33_w69, c0_n33_w70, c0_n33_w71, c0_n33_w72, c0_n33_w73, c0_n33_w74, c0_n33_w75, c0_n33_w76, c0_n33_w77, c0_n33_w78, c0_n33_w79, c0_n33_w80, c0_n33_w81, c0_n33_w82, c0_n33_w83, c0_n33_w84, c0_n33_w85, c0_n33_w86, c0_n33_w87, c0_n33_w88, c0_n33_w89, c0_n33_w90, c0_n33_w91, c0_n33_w92, c0_n33_w93, c0_n33_w94, c0_n33_w95, c0_n33_w96, c0_n33_w97, c0_n33_w98, c0_n33_w99, c0_n33_w100, c0_n33_w101, c0_n33_w102, c0_n33_w103, c0_n33_w104, c0_n33_w105, c0_n33_w106, c0_n33_w107, c0_n33_w108, c0_n33_w109, c0_n33_w110, c0_n33_w111, c0_n33_w112, c0_n33_w113, c0_n33_w114, c0_n33_w115, c0_n33_w116, c0_n33_w117, c0_n33_w118, c0_n33_w119, c0_n33_w120, c0_n33_w121, c0_n33_w122, c0_n33_w123, c0_n33_w124, c0_n33_w125, c0_n33_w126, c0_n33_w127, c0_n33_w128, c0_n33_w129, c0_n33_w130, c0_n33_w131, c0_n33_w132, c0_n33_w133, c0_n33_w134, c0_n33_w135, c0_n33_w136, c0_n33_w137, c0_n33_w138, c0_n33_w139, c0_n33_w140, c0_n33_w141, c0_n33_w142, c0_n33_w143, c0_n33_w144, c0_n33_w145, c0_n33_w146, c0_n33_w147, c0_n33_w148, c0_n33_w149, c0_n33_w150, c0_n33_w151, c0_n33_w152, c0_n33_w153, c0_n33_w154, c0_n33_w155, c0_n33_w156, c0_n33_w157, c0_n33_w158, c0_n33_w159, c0_n33_w160, c0_n33_w161, c0_n33_w162, c0_n33_w163, c0_n33_w164, c0_n33_w165, c0_n33_w166, c0_n33_w167, c0_n33_w168, c0_n33_w169, c0_n33_w170, c0_n33_w171, c0_n33_w172, c0_n33_w173, c0_n33_w174, c0_n33_w175, c0_n33_w176, c0_n33_w177, c0_n33_w178, c0_n33_w179, c0_n33_w180, c0_n33_w181, c0_n33_w182, c0_n33_w183, c0_n33_w184, c0_n33_w185, c0_n33_w186, c0_n33_w187, c0_n33_w188, c0_n33_w189, c0_n33_w190, c0_n33_w191, c0_n33_w192, c0_n33_w193, c0_n33_w194, c0_n33_w195, c0_n33_w196, c0_n33_w197, c0_n33_w198, c0_n33_w199, c0_n33_w200, c0_n34_w1, c0_n34_w2, c0_n34_w3, c0_n34_w4, c0_n34_w5, c0_n34_w6, c0_n34_w7, c0_n34_w8, c0_n34_w9, c0_n34_w10, c0_n34_w11, c0_n34_w12, c0_n34_w13, c0_n34_w14, c0_n34_w15, c0_n34_w16, c0_n34_w17, c0_n34_w18, c0_n34_w19, c0_n34_w20, c0_n34_w21, c0_n34_w22, c0_n34_w23, c0_n34_w24, c0_n34_w25, c0_n34_w26, c0_n34_w27, c0_n34_w28, c0_n34_w29, c0_n34_w30, c0_n34_w31, c0_n34_w32, c0_n34_w33, c0_n34_w34, c0_n34_w35, c0_n34_w36, c0_n34_w37, c0_n34_w38, c0_n34_w39, c0_n34_w40, c0_n34_w41, c0_n34_w42, c0_n34_w43, c0_n34_w44, c0_n34_w45, c0_n34_w46, c0_n34_w47, c0_n34_w48, c0_n34_w49, c0_n34_w50, c0_n34_w51, c0_n34_w52, c0_n34_w53, c0_n34_w54, c0_n34_w55, c0_n34_w56, c0_n34_w57, c0_n34_w58, c0_n34_w59, c0_n34_w60, c0_n34_w61, c0_n34_w62, c0_n34_w63, c0_n34_w64, c0_n34_w65, c0_n34_w66, c0_n34_w67, c0_n34_w68, c0_n34_w69, c0_n34_w70, c0_n34_w71, c0_n34_w72, c0_n34_w73, c0_n34_w74, c0_n34_w75, c0_n34_w76, c0_n34_w77, c0_n34_w78, c0_n34_w79, c0_n34_w80, c0_n34_w81, c0_n34_w82, c0_n34_w83, c0_n34_w84, c0_n34_w85, c0_n34_w86, c0_n34_w87, c0_n34_w88, c0_n34_w89, c0_n34_w90, c0_n34_w91, c0_n34_w92, c0_n34_w93, c0_n34_w94, c0_n34_w95, c0_n34_w96, c0_n34_w97, c0_n34_w98, c0_n34_w99, c0_n34_w100, c0_n34_w101, c0_n34_w102, c0_n34_w103, c0_n34_w104, c0_n34_w105, c0_n34_w106, c0_n34_w107, c0_n34_w108, c0_n34_w109, c0_n34_w110, c0_n34_w111, c0_n34_w112, c0_n34_w113, c0_n34_w114, c0_n34_w115, c0_n34_w116, c0_n34_w117, c0_n34_w118, c0_n34_w119, c0_n34_w120, c0_n34_w121, c0_n34_w122, c0_n34_w123, c0_n34_w124, c0_n34_w125, c0_n34_w126, c0_n34_w127, c0_n34_w128, c0_n34_w129, c0_n34_w130, c0_n34_w131, c0_n34_w132, c0_n34_w133, c0_n34_w134, c0_n34_w135, c0_n34_w136, c0_n34_w137, c0_n34_w138, c0_n34_w139, c0_n34_w140, c0_n34_w141, c0_n34_w142, c0_n34_w143, c0_n34_w144, c0_n34_w145, c0_n34_w146, c0_n34_w147, c0_n34_w148, c0_n34_w149, c0_n34_w150, c0_n34_w151, c0_n34_w152, c0_n34_w153, c0_n34_w154, c0_n34_w155, c0_n34_w156, c0_n34_w157, c0_n34_w158, c0_n34_w159, c0_n34_w160, c0_n34_w161, c0_n34_w162, c0_n34_w163, c0_n34_w164, c0_n34_w165, c0_n34_w166, c0_n34_w167, c0_n34_w168, c0_n34_w169, c0_n34_w170, c0_n34_w171, c0_n34_w172, c0_n34_w173, c0_n34_w174, c0_n34_w175, c0_n34_w176, c0_n34_w177, c0_n34_w178, c0_n34_w179, c0_n34_w180, c0_n34_w181, c0_n34_w182, c0_n34_w183, c0_n34_w184, c0_n34_w185, c0_n34_w186, c0_n34_w187, c0_n34_w188, c0_n34_w189, c0_n34_w190, c0_n34_w191, c0_n34_w192, c0_n34_w193, c0_n34_w194, c0_n34_w195, c0_n34_w196, c0_n34_w197, c0_n34_w198, c0_n34_w199, c0_n34_w200, c0_n35_w1, c0_n35_w2, c0_n35_w3, c0_n35_w4, c0_n35_w5, c0_n35_w6, c0_n35_w7, c0_n35_w8, c0_n35_w9, c0_n35_w10, c0_n35_w11, c0_n35_w12, c0_n35_w13, c0_n35_w14, c0_n35_w15, c0_n35_w16, c0_n35_w17, c0_n35_w18, c0_n35_w19, c0_n35_w20, c0_n35_w21, c0_n35_w22, c0_n35_w23, c0_n35_w24, c0_n35_w25, c0_n35_w26, c0_n35_w27, c0_n35_w28, c0_n35_w29, c0_n35_w30, c0_n35_w31, c0_n35_w32, c0_n35_w33, c0_n35_w34, c0_n35_w35, c0_n35_w36, c0_n35_w37, c0_n35_w38, c0_n35_w39, c0_n35_w40, c0_n35_w41, c0_n35_w42, c0_n35_w43, c0_n35_w44, c0_n35_w45, c0_n35_w46, c0_n35_w47, c0_n35_w48, c0_n35_w49, c0_n35_w50, c0_n35_w51, c0_n35_w52, c0_n35_w53, c0_n35_w54, c0_n35_w55, c0_n35_w56, c0_n35_w57, c0_n35_w58, c0_n35_w59, c0_n35_w60, c0_n35_w61, c0_n35_w62, c0_n35_w63, c0_n35_w64, c0_n35_w65, c0_n35_w66, c0_n35_w67, c0_n35_w68, c0_n35_w69, c0_n35_w70, c0_n35_w71, c0_n35_w72, c0_n35_w73, c0_n35_w74, c0_n35_w75, c0_n35_w76, c0_n35_w77, c0_n35_w78, c0_n35_w79, c0_n35_w80, c0_n35_w81, c0_n35_w82, c0_n35_w83, c0_n35_w84, c0_n35_w85, c0_n35_w86, c0_n35_w87, c0_n35_w88, c0_n35_w89, c0_n35_w90, c0_n35_w91, c0_n35_w92, c0_n35_w93, c0_n35_w94, c0_n35_w95, c0_n35_w96, c0_n35_w97, c0_n35_w98, c0_n35_w99, c0_n35_w100, c0_n35_w101, c0_n35_w102, c0_n35_w103, c0_n35_w104, c0_n35_w105, c0_n35_w106, c0_n35_w107, c0_n35_w108, c0_n35_w109, c0_n35_w110, c0_n35_w111, c0_n35_w112, c0_n35_w113, c0_n35_w114, c0_n35_w115, c0_n35_w116, c0_n35_w117, c0_n35_w118, c0_n35_w119, c0_n35_w120, c0_n35_w121, c0_n35_w122, c0_n35_w123, c0_n35_w124, c0_n35_w125, c0_n35_w126, c0_n35_w127, c0_n35_w128, c0_n35_w129, c0_n35_w130, c0_n35_w131, c0_n35_w132, c0_n35_w133, c0_n35_w134, c0_n35_w135, c0_n35_w136, c0_n35_w137, c0_n35_w138, c0_n35_w139, c0_n35_w140, c0_n35_w141, c0_n35_w142, c0_n35_w143, c0_n35_w144, c0_n35_w145, c0_n35_w146, c0_n35_w147, c0_n35_w148, c0_n35_w149, c0_n35_w150, c0_n35_w151, c0_n35_w152, c0_n35_w153, c0_n35_w154, c0_n35_w155, c0_n35_w156, c0_n35_w157, c0_n35_w158, c0_n35_w159, c0_n35_w160, c0_n35_w161, c0_n35_w162, c0_n35_w163, c0_n35_w164, c0_n35_w165, c0_n35_w166, c0_n35_w167, c0_n35_w168, c0_n35_w169, c0_n35_w170, c0_n35_w171, c0_n35_w172, c0_n35_w173, c0_n35_w174, c0_n35_w175, c0_n35_w176, c0_n35_w177, c0_n35_w178, c0_n35_w179, c0_n35_w180, c0_n35_w181, c0_n35_w182, c0_n35_w183, c0_n35_w184, c0_n35_w185, c0_n35_w186, c0_n35_w187, c0_n35_w188, c0_n35_w189, c0_n35_w190, c0_n35_w191, c0_n35_w192, c0_n35_w193, c0_n35_w194, c0_n35_w195, c0_n35_w196, c0_n35_w197, c0_n35_w198, c0_n35_w199, c0_n35_w200, c0_n36_w1, c0_n36_w2, c0_n36_w3, c0_n36_w4, c0_n36_w5, c0_n36_w6, c0_n36_w7, c0_n36_w8, c0_n36_w9, c0_n36_w10, c0_n36_w11, c0_n36_w12, c0_n36_w13, c0_n36_w14, c0_n36_w15, c0_n36_w16, c0_n36_w17, c0_n36_w18, c0_n36_w19, c0_n36_w20, c0_n36_w21, c0_n36_w22, c0_n36_w23, c0_n36_w24, c0_n36_w25, c0_n36_w26, c0_n36_w27, c0_n36_w28, c0_n36_w29, c0_n36_w30, c0_n36_w31, c0_n36_w32, c0_n36_w33, c0_n36_w34, c0_n36_w35, c0_n36_w36, c0_n36_w37, c0_n36_w38, c0_n36_w39, c0_n36_w40, c0_n36_w41, c0_n36_w42, c0_n36_w43, c0_n36_w44, c0_n36_w45, c0_n36_w46, c0_n36_w47, c0_n36_w48, c0_n36_w49, c0_n36_w50, c0_n36_w51, c0_n36_w52, c0_n36_w53, c0_n36_w54, c0_n36_w55, c0_n36_w56, c0_n36_w57, c0_n36_w58, c0_n36_w59, c0_n36_w60, c0_n36_w61, c0_n36_w62, c0_n36_w63, c0_n36_w64, c0_n36_w65, c0_n36_w66, c0_n36_w67, c0_n36_w68, c0_n36_w69, c0_n36_w70, c0_n36_w71, c0_n36_w72, c0_n36_w73, c0_n36_w74, c0_n36_w75, c0_n36_w76, c0_n36_w77, c0_n36_w78, c0_n36_w79, c0_n36_w80, c0_n36_w81, c0_n36_w82, c0_n36_w83, c0_n36_w84, c0_n36_w85, c0_n36_w86, c0_n36_w87, c0_n36_w88, c0_n36_w89, c0_n36_w90, c0_n36_w91, c0_n36_w92, c0_n36_w93, c0_n36_w94, c0_n36_w95, c0_n36_w96, c0_n36_w97, c0_n36_w98, c0_n36_w99, c0_n36_w100, c0_n36_w101, c0_n36_w102, c0_n36_w103, c0_n36_w104, c0_n36_w105, c0_n36_w106, c0_n36_w107, c0_n36_w108, c0_n36_w109, c0_n36_w110, c0_n36_w111, c0_n36_w112, c0_n36_w113, c0_n36_w114, c0_n36_w115, c0_n36_w116, c0_n36_w117, c0_n36_w118, c0_n36_w119, c0_n36_w120, c0_n36_w121, c0_n36_w122, c0_n36_w123, c0_n36_w124, c0_n36_w125, c0_n36_w126, c0_n36_w127, c0_n36_w128, c0_n36_w129, c0_n36_w130, c0_n36_w131, c0_n36_w132, c0_n36_w133, c0_n36_w134, c0_n36_w135, c0_n36_w136, c0_n36_w137, c0_n36_w138, c0_n36_w139, c0_n36_w140, c0_n36_w141, c0_n36_w142, c0_n36_w143, c0_n36_w144, c0_n36_w145, c0_n36_w146, c0_n36_w147, c0_n36_w148, c0_n36_w149, c0_n36_w150, c0_n36_w151, c0_n36_w152, c0_n36_w153, c0_n36_w154, c0_n36_w155, c0_n36_w156, c0_n36_w157, c0_n36_w158, c0_n36_w159, c0_n36_w160, c0_n36_w161, c0_n36_w162, c0_n36_w163, c0_n36_w164, c0_n36_w165, c0_n36_w166, c0_n36_w167, c0_n36_w168, c0_n36_w169, c0_n36_w170, c0_n36_w171, c0_n36_w172, c0_n36_w173, c0_n36_w174, c0_n36_w175, c0_n36_w176, c0_n36_w177, c0_n36_w178, c0_n36_w179, c0_n36_w180, c0_n36_w181, c0_n36_w182, c0_n36_w183, c0_n36_w184, c0_n36_w185, c0_n36_w186, c0_n36_w187, c0_n36_w188, c0_n36_w189, c0_n36_w190, c0_n36_w191, c0_n36_w192, c0_n36_w193, c0_n36_w194, c0_n36_w195, c0_n36_w196, c0_n36_w197, c0_n36_w198, c0_n36_w199, c0_n36_w200, c0_n37_w1, c0_n37_w2, c0_n37_w3, c0_n37_w4, c0_n37_w5, c0_n37_w6, c0_n37_w7, c0_n37_w8, c0_n37_w9, c0_n37_w10, c0_n37_w11, c0_n37_w12, c0_n37_w13, c0_n37_w14, c0_n37_w15, c0_n37_w16, c0_n37_w17, c0_n37_w18, c0_n37_w19, c0_n37_w20, c0_n37_w21, c0_n37_w22, c0_n37_w23, c0_n37_w24, c0_n37_w25, c0_n37_w26, c0_n37_w27, c0_n37_w28, c0_n37_w29, c0_n37_w30, c0_n37_w31, c0_n37_w32, c0_n37_w33, c0_n37_w34, c0_n37_w35, c0_n37_w36, c0_n37_w37, c0_n37_w38, c0_n37_w39, c0_n37_w40, c0_n37_w41, c0_n37_w42, c0_n37_w43, c0_n37_w44, c0_n37_w45, c0_n37_w46, c0_n37_w47, c0_n37_w48, c0_n37_w49, c0_n37_w50, c0_n37_w51, c0_n37_w52, c0_n37_w53, c0_n37_w54, c0_n37_w55, c0_n37_w56, c0_n37_w57, c0_n37_w58, c0_n37_w59, c0_n37_w60, c0_n37_w61, c0_n37_w62, c0_n37_w63, c0_n37_w64, c0_n37_w65, c0_n37_w66, c0_n37_w67, c0_n37_w68, c0_n37_w69, c0_n37_w70, c0_n37_w71, c0_n37_w72, c0_n37_w73, c0_n37_w74, c0_n37_w75, c0_n37_w76, c0_n37_w77, c0_n37_w78, c0_n37_w79, c0_n37_w80, c0_n37_w81, c0_n37_w82, c0_n37_w83, c0_n37_w84, c0_n37_w85, c0_n37_w86, c0_n37_w87, c0_n37_w88, c0_n37_w89, c0_n37_w90, c0_n37_w91, c0_n37_w92, c0_n37_w93, c0_n37_w94, c0_n37_w95, c0_n37_w96, c0_n37_w97, c0_n37_w98, c0_n37_w99, c0_n37_w100, c0_n37_w101, c0_n37_w102, c0_n37_w103, c0_n37_w104, c0_n37_w105, c0_n37_w106, c0_n37_w107, c0_n37_w108, c0_n37_w109, c0_n37_w110, c0_n37_w111, c0_n37_w112, c0_n37_w113, c0_n37_w114, c0_n37_w115, c0_n37_w116, c0_n37_w117, c0_n37_w118, c0_n37_w119, c0_n37_w120, c0_n37_w121, c0_n37_w122, c0_n37_w123, c0_n37_w124, c0_n37_w125, c0_n37_w126, c0_n37_w127, c0_n37_w128, c0_n37_w129, c0_n37_w130, c0_n37_w131, c0_n37_w132, c0_n37_w133, c0_n37_w134, c0_n37_w135, c0_n37_w136, c0_n37_w137, c0_n37_w138, c0_n37_w139, c0_n37_w140, c0_n37_w141, c0_n37_w142, c0_n37_w143, c0_n37_w144, c0_n37_w145, c0_n37_w146, c0_n37_w147, c0_n37_w148, c0_n37_w149, c0_n37_w150, c0_n37_w151, c0_n37_w152, c0_n37_w153, c0_n37_w154, c0_n37_w155, c0_n37_w156, c0_n37_w157, c0_n37_w158, c0_n37_w159, c0_n37_w160, c0_n37_w161, c0_n37_w162, c0_n37_w163, c0_n37_w164, c0_n37_w165, c0_n37_w166, c0_n37_w167, c0_n37_w168, c0_n37_w169, c0_n37_w170, c0_n37_w171, c0_n37_w172, c0_n37_w173, c0_n37_w174, c0_n37_w175, c0_n37_w176, c0_n37_w177, c0_n37_w178, c0_n37_w179, c0_n37_w180, c0_n37_w181, c0_n37_w182, c0_n37_w183, c0_n37_w184, c0_n37_w185, c0_n37_w186, c0_n37_w187, c0_n37_w188, c0_n37_w189, c0_n37_w190, c0_n37_w191, c0_n37_w192, c0_n37_w193, c0_n37_w194, c0_n37_w195, c0_n37_w196, c0_n37_w197, c0_n37_w198, c0_n37_w199, c0_n37_w200, c0_n38_w1, c0_n38_w2, c0_n38_w3, c0_n38_w4, c0_n38_w5, c0_n38_w6, c0_n38_w7, c0_n38_w8, c0_n38_w9, c0_n38_w10, c0_n38_w11, c0_n38_w12, c0_n38_w13, c0_n38_w14, c0_n38_w15, c0_n38_w16, c0_n38_w17, c0_n38_w18, c0_n38_w19, c0_n38_w20, c0_n38_w21, c0_n38_w22, c0_n38_w23, c0_n38_w24, c0_n38_w25, c0_n38_w26, c0_n38_w27, c0_n38_w28, c0_n38_w29, c0_n38_w30, c0_n38_w31, c0_n38_w32, c0_n38_w33, c0_n38_w34, c0_n38_w35, c0_n38_w36, c0_n38_w37, c0_n38_w38, c0_n38_w39, c0_n38_w40, c0_n38_w41, c0_n38_w42, c0_n38_w43, c0_n38_w44, c0_n38_w45, c0_n38_w46, c0_n38_w47, c0_n38_w48, c0_n38_w49, c0_n38_w50, c0_n38_w51, c0_n38_w52, c0_n38_w53, c0_n38_w54, c0_n38_w55, c0_n38_w56, c0_n38_w57, c0_n38_w58, c0_n38_w59, c0_n38_w60, c0_n38_w61, c0_n38_w62, c0_n38_w63, c0_n38_w64, c0_n38_w65, c0_n38_w66, c0_n38_w67, c0_n38_w68, c0_n38_w69, c0_n38_w70, c0_n38_w71, c0_n38_w72, c0_n38_w73, c0_n38_w74, c0_n38_w75, c0_n38_w76, c0_n38_w77, c0_n38_w78, c0_n38_w79, c0_n38_w80, c0_n38_w81, c0_n38_w82, c0_n38_w83, c0_n38_w84, c0_n38_w85, c0_n38_w86, c0_n38_w87, c0_n38_w88, c0_n38_w89, c0_n38_w90, c0_n38_w91, c0_n38_w92, c0_n38_w93, c0_n38_w94, c0_n38_w95, c0_n38_w96, c0_n38_w97, c0_n38_w98, c0_n38_w99, c0_n38_w100, c0_n38_w101, c0_n38_w102, c0_n38_w103, c0_n38_w104, c0_n38_w105, c0_n38_w106, c0_n38_w107, c0_n38_w108, c0_n38_w109, c0_n38_w110, c0_n38_w111, c0_n38_w112, c0_n38_w113, c0_n38_w114, c0_n38_w115, c0_n38_w116, c0_n38_w117, c0_n38_w118, c0_n38_w119, c0_n38_w120, c0_n38_w121, c0_n38_w122, c0_n38_w123, c0_n38_w124, c0_n38_w125, c0_n38_w126, c0_n38_w127, c0_n38_w128, c0_n38_w129, c0_n38_w130, c0_n38_w131, c0_n38_w132, c0_n38_w133, c0_n38_w134, c0_n38_w135, c0_n38_w136, c0_n38_w137, c0_n38_w138, c0_n38_w139, c0_n38_w140, c0_n38_w141, c0_n38_w142, c0_n38_w143, c0_n38_w144, c0_n38_w145, c0_n38_w146, c0_n38_w147, c0_n38_w148, c0_n38_w149, c0_n38_w150, c0_n38_w151, c0_n38_w152, c0_n38_w153, c0_n38_w154, c0_n38_w155, c0_n38_w156, c0_n38_w157, c0_n38_w158, c0_n38_w159, c0_n38_w160, c0_n38_w161, c0_n38_w162, c0_n38_w163, c0_n38_w164, c0_n38_w165, c0_n38_w166, c0_n38_w167, c0_n38_w168, c0_n38_w169, c0_n38_w170, c0_n38_w171, c0_n38_w172, c0_n38_w173, c0_n38_w174, c0_n38_w175, c0_n38_w176, c0_n38_w177, c0_n38_w178, c0_n38_w179, c0_n38_w180, c0_n38_w181, c0_n38_w182, c0_n38_w183, c0_n38_w184, c0_n38_w185, c0_n38_w186, c0_n38_w187, c0_n38_w188, c0_n38_w189, c0_n38_w190, c0_n38_w191, c0_n38_w192, c0_n38_w193, c0_n38_w194, c0_n38_w195, c0_n38_w196, c0_n38_w197, c0_n38_w198, c0_n38_w199, c0_n38_w200, c0_n39_w1, c0_n39_w2, c0_n39_w3, c0_n39_w4, c0_n39_w5, c0_n39_w6, c0_n39_w7, c0_n39_w8, c0_n39_w9, c0_n39_w10, c0_n39_w11, c0_n39_w12, c0_n39_w13, c0_n39_w14, c0_n39_w15, c0_n39_w16, c0_n39_w17, c0_n39_w18, c0_n39_w19, c0_n39_w20, c0_n39_w21, c0_n39_w22, c0_n39_w23, c0_n39_w24, c0_n39_w25, c0_n39_w26, c0_n39_w27, c0_n39_w28, c0_n39_w29, c0_n39_w30, c0_n39_w31, c0_n39_w32, c0_n39_w33, c0_n39_w34, c0_n39_w35, c0_n39_w36, c0_n39_w37, c0_n39_w38, c0_n39_w39, c0_n39_w40, c0_n39_w41, c0_n39_w42, c0_n39_w43, c0_n39_w44, c0_n39_w45, c0_n39_w46, c0_n39_w47, c0_n39_w48, c0_n39_w49, c0_n39_w50, c0_n39_w51, c0_n39_w52, c0_n39_w53, c0_n39_w54, c0_n39_w55, c0_n39_w56, c0_n39_w57, c0_n39_w58, c0_n39_w59, c0_n39_w60, c0_n39_w61, c0_n39_w62, c0_n39_w63, c0_n39_w64, c0_n39_w65, c0_n39_w66, c0_n39_w67, c0_n39_w68, c0_n39_w69, c0_n39_w70, c0_n39_w71, c0_n39_w72, c0_n39_w73, c0_n39_w74, c0_n39_w75, c0_n39_w76, c0_n39_w77, c0_n39_w78, c0_n39_w79, c0_n39_w80, c0_n39_w81, c0_n39_w82, c0_n39_w83, c0_n39_w84, c0_n39_w85, c0_n39_w86, c0_n39_w87, c0_n39_w88, c0_n39_w89, c0_n39_w90, c0_n39_w91, c0_n39_w92, c0_n39_w93, c0_n39_w94, c0_n39_w95, c0_n39_w96, c0_n39_w97, c0_n39_w98, c0_n39_w99, c0_n39_w100, c0_n39_w101, c0_n39_w102, c0_n39_w103, c0_n39_w104, c0_n39_w105, c0_n39_w106, c0_n39_w107, c0_n39_w108, c0_n39_w109, c0_n39_w110, c0_n39_w111, c0_n39_w112, c0_n39_w113, c0_n39_w114, c0_n39_w115, c0_n39_w116, c0_n39_w117, c0_n39_w118, c0_n39_w119, c0_n39_w120, c0_n39_w121, c0_n39_w122, c0_n39_w123, c0_n39_w124, c0_n39_w125, c0_n39_w126, c0_n39_w127, c0_n39_w128, c0_n39_w129, c0_n39_w130, c0_n39_w131, c0_n39_w132, c0_n39_w133, c0_n39_w134, c0_n39_w135, c0_n39_w136, c0_n39_w137, c0_n39_w138, c0_n39_w139, c0_n39_w140, c0_n39_w141, c0_n39_w142, c0_n39_w143, c0_n39_w144, c0_n39_w145, c0_n39_w146, c0_n39_w147, c0_n39_w148, c0_n39_w149, c0_n39_w150, c0_n39_w151, c0_n39_w152, c0_n39_w153, c0_n39_w154, c0_n39_w155, c0_n39_w156, c0_n39_w157, c0_n39_w158, c0_n39_w159, c0_n39_w160, c0_n39_w161, c0_n39_w162, c0_n39_w163, c0_n39_w164, c0_n39_w165, c0_n39_w166, c0_n39_w167, c0_n39_w168, c0_n39_w169, c0_n39_w170, c0_n39_w171, c0_n39_w172, c0_n39_w173, c0_n39_w174, c0_n39_w175, c0_n39_w176, c0_n39_w177, c0_n39_w178, c0_n39_w179, c0_n39_w180, c0_n39_w181, c0_n39_w182, c0_n39_w183, c0_n39_w184, c0_n39_w185, c0_n39_w186, c0_n39_w187, c0_n39_w188, c0_n39_w189, c0_n39_w190, c0_n39_w191, c0_n39_w192, c0_n39_w193, c0_n39_w194, c0_n39_w195, c0_n39_w196, c0_n39_w197, c0_n39_w198, c0_n39_w199, c0_n39_w200, c0_n40_w1, c0_n40_w2, c0_n40_w3, c0_n40_w4, c0_n40_w5, c0_n40_w6, c0_n40_w7, c0_n40_w8, c0_n40_w9, c0_n40_w10, c0_n40_w11, c0_n40_w12, c0_n40_w13, c0_n40_w14, c0_n40_w15, c0_n40_w16, c0_n40_w17, c0_n40_w18, c0_n40_w19, c0_n40_w20, c0_n40_w21, c0_n40_w22, c0_n40_w23, c0_n40_w24, c0_n40_w25, c0_n40_w26, c0_n40_w27, c0_n40_w28, c0_n40_w29, c0_n40_w30, c0_n40_w31, c0_n40_w32, c0_n40_w33, c0_n40_w34, c0_n40_w35, c0_n40_w36, c0_n40_w37, c0_n40_w38, c0_n40_w39, c0_n40_w40, c0_n40_w41, c0_n40_w42, c0_n40_w43, c0_n40_w44, c0_n40_w45, c0_n40_w46, c0_n40_w47, c0_n40_w48, c0_n40_w49, c0_n40_w50, c0_n40_w51, c0_n40_w52, c0_n40_w53, c0_n40_w54, c0_n40_w55, c0_n40_w56, c0_n40_w57, c0_n40_w58, c0_n40_w59, c0_n40_w60, c0_n40_w61, c0_n40_w62, c0_n40_w63, c0_n40_w64, c0_n40_w65, c0_n40_w66, c0_n40_w67, c0_n40_w68, c0_n40_w69, c0_n40_w70, c0_n40_w71, c0_n40_w72, c0_n40_w73, c0_n40_w74, c0_n40_w75, c0_n40_w76, c0_n40_w77, c0_n40_w78, c0_n40_w79, c0_n40_w80, c0_n40_w81, c0_n40_w82, c0_n40_w83, c0_n40_w84, c0_n40_w85, c0_n40_w86, c0_n40_w87, c0_n40_w88, c0_n40_w89, c0_n40_w90, c0_n40_w91, c0_n40_w92, c0_n40_w93, c0_n40_w94, c0_n40_w95, c0_n40_w96, c0_n40_w97, c0_n40_w98, c0_n40_w99, c0_n40_w100, c0_n40_w101, c0_n40_w102, c0_n40_w103, c0_n40_w104, c0_n40_w105, c0_n40_w106, c0_n40_w107, c0_n40_w108, c0_n40_w109, c0_n40_w110, c0_n40_w111, c0_n40_w112, c0_n40_w113, c0_n40_w114, c0_n40_w115, c0_n40_w116, c0_n40_w117, c0_n40_w118, c0_n40_w119, c0_n40_w120, c0_n40_w121, c0_n40_w122, c0_n40_w123, c0_n40_w124, c0_n40_w125, c0_n40_w126, c0_n40_w127, c0_n40_w128, c0_n40_w129, c0_n40_w130, c0_n40_w131, c0_n40_w132, c0_n40_w133, c0_n40_w134, c0_n40_w135, c0_n40_w136, c0_n40_w137, c0_n40_w138, c0_n40_w139, c0_n40_w140, c0_n40_w141, c0_n40_w142, c0_n40_w143, c0_n40_w144, c0_n40_w145, c0_n40_w146, c0_n40_w147, c0_n40_w148, c0_n40_w149, c0_n40_w150, c0_n40_w151, c0_n40_w152, c0_n40_w153, c0_n40_w154, c0_n40_w155, c0_n40_w156, c0_n40_w157, c0_n40_w158, c0_n40_w159, c0_n40_w160, c0_n40_w161, c0_n40_w162, c0_n40_w163, c0_n40_w164, c0_n40_w165, c0_n40_w166, c0_n40_w167, c0_n40_w168, c0_n40_w169, c0_n40_w170, c0_n40_w171, c0_n40_w172, c0_n40_w173, c0_n40_w174, c0_n40_w175, c0_n40_w176, c0_n40_w177, c0_n40_w178, c0_n40_w179, c0_n40_w180, c0_n40_w181, c0_n40_w182, c0_n40_w183, c0_n40_w184, c0_n40_w185, c0_n40_w186, c0_n40_w187, c0_n40_w188, c0_n40_w189, c0_n40_w190, c0_n40_w191, c0_n40_w192, c0_n40_w193, c0_n40_w194, c0_n40_w195, c0_n40_w196, c0_n40_w197, c0_n40_w198, c0_n40_w199, c0_n40_w200, c0_n41_w1, c0_n41_w2, c0_n41_w3, c0_n41_w4, c0_n41_w5, c0_n41_w6, c0_n41_w7, c0_n41_w8, c0_n41_w9, c0_n41_w10, c0_n41_w11, c0_n41_w12, c0_n41_w13, c0_n41_w14, c0_n41_w15, c0_n41_w16, c0_n41_w17, c0_n41_w18, c0_n41_w19, c0_n41_w20, c0_n41_w21, c0_n41_w22, c0_n41_w23, c0_n41_w24, c0_n41_w25, c0_n41_w26, c0_n41_w27, c0_n41_w28, c0_n41_w29, c0_n41_w30, c0_n41_w31, c0_n41_w32, c0_n41_w33, c0_n41_w34, c0_n41_w35, c0_n41_w36, c0_n41_w37, c0_n41_w38, c0_n41_w39, c0_n41_w40, c0_n41_w41, c0_n41_w42, c0_n41_w43, c0_n41_w44, c0_n41_w45, c0_n41_w46, c0_n41_w47, c0_n41_w48, c0_n41_w49, c0_n41_w50, c0_n41_w51, c0_n41_w52, c0_n41_w53, c0_n41_w54, c0_n41_w55, c0_n41_w56, c0_n41_w57, c0_n41_w58, c0_n41_w59, c0_n41_w60, c0_n41_w61, c0_n41_w62, c0_n41_w63, c0_n41_w64, c0_n41_w65, c0_n41_w66, c0_n41_w67, c0_n41_w68, c0_n41_w69, c0_n41_w70, c0_n41_w71, c0_n41_w72, c0_n41_w73, c0_n41_w74, c0_n41_w75, c0_n41_w76, c0_n41_w77, c0_n41_w78, c0_n41_w79, c0_n41_w80, c0_n41_w81, c0_n41_w82, c0_n41_w83, c0_n41_w84, c0_n41_w85, c0_n41_w86, c0_n41_w87, c0_n41_w88, c0_n41_w89, c0_n41_w90, c0_n41_w91, c0_n41_w92, c0_n41_w93, c0_n41_w94, c0_n41_w95, c0_n41_w96, c0_n41_w97, c0_n41_w98, c0_n41_w99, c0_n41_w100, c0_n41_w101, c0_n41_w102, c0_n41_w103, c0_n41_w104, c0_n41_w105, c0_n41_w106, c0_n41_w107, c0_n41_w108, c0_n41_w109, c0_n41_w110, c0_n41_w111, c0_n41_w112, c0_n41_w113, c0_n41_w114, c0_n41_w115, c0_n41_w116, c0_n41_w117, c0_n41_w118, c0_n41_w119, c0_n41_w120, c0_n41_w121, c0_n41_w122, c0_n41_w123, c0_n41_w124, c0_n41_w125, c0_n41_w126, c0_n41_w127, c0_n41_w128, c0_n41_w129, c0_n41_w130, c0_n41_w131, c0_n41_w132, c0_n41_w133, c0_n41_w134, c0_n41_w135, c0_n41_w136, c0_n41_w137, c0_n41_w138, c0_n41_w139, c0_n41_w140, c0_n41_w141, c0_n41_w142, c0_n41_w143, c0_n41_w144, c0_n41_w145, c0_n41_w146, c0_n41_w147, c0_n41_w148, c0_n41_w149, c0_n41_w150, c0_n41_w151, c0_n41_w152, c0_n41_w153, c0_n41_w154, c0_n41_w155, c0_n41_w156, c0_n41_w157, c0_n41_w158, c0_n41_w159, c0_n41_w160, c0_n41_w161, c0_n41_w162, c0_n41_w163, c0_n41_w164, c0_n41_w165, c0_n41_w166, c0_n41_w167, c0_n41_w168, c0_n41_w169, c0_n41_w170, c0_n41_w171, c0_n41_w172, c0_n41_w173, c0_n41_w174, c0_n41_w175, c0_n41_w176, c0_n41_w177, c0_n41_w178, c0_n41_w179, c0_n41_w180, c0_n41_w181, c0_n41_w182, c0_n41_w183, c0_n41_w184, c0_n41_w185, c0_n41_w186, c0_n41_w187, c0_n41_w188, c0_n41_w189, c0_n41_w190, c0_n41_w191, c0_n41_w192, c0_n41_w193, c0_n41_w194, c0_n41_w195, c0_n41_w196, c0_n41_w197, c0_n41_w198, c0_n41_w199, c0_n41_w200, c0_n42_w1, c0_n42_w2, c0_n42_w3, c0_n42_w4, c0_n42_w5, c0_n42_w6, c0_n42_w7, c0_n42_w8, c0_n42_w9, c0_n42_w10, c0_n42_w11, c0_n42_w12, c0_n42_w13, c0_n42_w14, c0_n42_w15, c0_n42_w16, c0_n42_w17, c0_n42_w18, c0_n42_w19, c0_n42_w20, c0_n42_w21, c0_n42_w22, c0_n42_w23, c0_n42_w24, c0_n42_w25, c0_n42_w26, c0_n42_w27, c0_n42_w28, c0_n42_w29, c0_n42_w30, c0_n42_w31, c0_n42_w32, c0_n42_w33, c0_n42_w34, c0_n42_w35, c0_n42_w36, c0_n42_w37, c0_n42_w38, c0_n42_w39, c0_n42_w40, c0_n42_w41, c0_n42_w42, c0_n42_w43, c0_n42_w44, c0_n42_w45, c0_n42_w46, c0_n42_w47, c0_n42_w48, c0_n42_w49, c0_n42_w50, c0_n42_w51, c0_n42_w52, c0_n42_w53, c0_n42_w54, c0_n42_w55, c0_n42_w56, c0_n42_w57, c0_n42_w58, c0_n42_w59, c0_n42_w60, c0_n42_w61, c0_n42_w62, c0_n42_w63, c0_n42_w64, c0_n42_w65, c0_n42_w66, c0_n42_w67, c0_n42_w68, c0_n42_w69, c0_n42_w70, c0_n42_w71, c0_n42_w72, c0_n42_w73, c0_n42_w74, c0_n42_w75, c0_n42_w76, c0_n42_w77, c0_n42_w78, c0_n42_w79, c0_n42_w80, c0_n42_w81, c0_n42_w82, c0_n42_w83, c0_n42_w84, c0_n42_w85, c0_n42_w86, c0_n42_w87, c0_n42_w88, c0_n42_w89, c0_n42_w90, c0_n42_w91, c0_n42_w92, c0_n42_w93, c0_n42_w94, c0_n42_w95, c0_n42_w96, c0_n42_w97, c0_n42_w98, c0_n42_w99, c0_n42_w100, c0_n42_w101, c0_n42_w102, c0_n42_w103, c0_n42_w104, c0_n42_w105, c0_n42_w106, c0_n42_w107, c0_n42_w108, c0_n42_w109, c0_n42_w110, c0_n42_w111, c0_n42_w112, c0_n42_w113, c0_n42_w114, c0_n42_w115, c0_n42_w116, c0_n42_w117, c0_n42_w118, c0_n42_w119, c0_n42_w120, c0_n42_w121, c0_n42_w122, c0_n42_w123, c0_n42_w124, c0_n42_w125, c0_n42_w126, c0_n42_w127, c0_n42_w128, c0_n42_w129, c0_n42_w130, c0_n42_w131, c0_n42_w132, c0_n42_w133, c0_n42_w134, c0_n42_w135, c0_n42_w136, c0_n42_w137, c0_n42_w138, c0_n42_w139, c0_n42_w140, c0_n42_w141, c0_n42_w142, c0_n42_w143, c0_n42_w144, c0_n42_w145, c0_n42_w146, c0_n42_w147, c0_n42_w148, c0_n42_w149, c0_n42_w150, c0_n42_w151, c0_n42_w152, c0_n42_w153, c0_n42_w154, c0_n42_w155, c0_n42_w156, c0_n42_w157, c0_n42_w158, c0_n42_w159, c0_n42_w160, c0_n42_w161, c0_n42_w162, c0_n42_w163, c0_n42_w164, c0_n42_w165, c0_n42_w166, c0_n42_w167, c0_n42_w168, c0_n42_w169, c0_n42_w170, c0_n42_w171, c0_n42_w172, c0_n42_w173, c0_n42_w174, c0_n42_w175, c0_n42_w176, c0_n42_w177, c0_n42_w178, c0_n42_w179, c0_n42_w180, c0_n42_w181, c0_n42_w182, c0_n42_w183, c0_n42_w184, c0_n42_w185, c0_n42_w186, c0_n42_w187, c0_n42_w188, c0_n42_w189, c0_n42_w190, c0_n42_w191, c0_n42_w192, c0_n42_w193, c0_n42_w194, c0_n42_w195, c0_n42_w196, c0_n42_w197, c0_n42_w198, c0_n42_w199, c0_n42_w200, c0_n43_w1, c0_n43_w2, c0_n43_w3, c0_n43_w4, c0_n43_w5, c0_n43_w6, c0_n43_w7, c0_n43_w8, c0_n43_w9, c0_n43_w10, c0_n43_w11, c0_n43_w12, c0_n43_w13, c0_n43_w14, c0_n43_w15, c0_n43_w16, c0_n43_w17, c0_n43_w18, c0_n43_w19, c0_n43_w20, c0_n43_w21, c0_n43_w22, c0_n43_w23, c0_n43_w24, c0_n43_w25, c0_n43_w26, c0_n43_w27, c0_n43_w28, c0_n43_w29, c0_n43_w30, c0_n43_w31, c0_n43_w32, c0_n43_w33, c0_n43_w34, c0_n43_w35, c0_n43_w36, c0_n43_w37, c0_n43_w38, c0_n43_w39, c0_n43_w40, c0_n43_w41, c0_n43_w42, c0_n43_w43, c0_n43_w44, c0_n43_w45, c0_n43_w46, c0_n43_w47, c0_n43_w48, c0_n43_w49, c0_n43_w50, c0_n43_w51, c0_n43_w52, c0_n43_w53, c0_n43_w54, c0_n43_w55, c0_n43_w56, c0_n43_w57, c0_n43_w58, c0_n43_w59, c0_n43_w60, c0_n43_w61, c0_n43_w62, c0_n43_w63, c0_n43_w64, c0_n43_w65, c0_n43_w66, c0_n43_w67, c0_n43_w68, c0_n43_w69, c0_n43_w70, c0_n43_w71, c0_n43_w72, c0_n43_w73, c0_n43_w74, c0_n43_w75, c0_n43_w76, c0_n43_w77, c0_n43_w78, c0_n43_w79, c0_n43_w80, c0_n43_w81, c0_n43_w82, c0_n43_w83, c0_n43_w84, c0_n43_w85, c0_n43_w86, c0_n43_w87, c0_n43_w88, c0_n43_w89, c0_n43_w90, c0_n43_w91, c0_n43_w92, c0_n43_w93, c0_n43_w94, c0_n43_w95, c0_n43_w96, c0_n43_w97, c0_n43_w98, c0_n43_w99, c0_n43_w100, c0_n43_w101, c0_n43_w102, c0_n43_w103, c0_n43_w104, c0_n43_w105, c0_n43_w106, c0_n43_w107, c0_n43_w108, c0_n43_w109, c0_n43_w110, c0_n43_w111, c0_n43_w112, c0_n43_w113, c0_n43_w114, c0_n43_w115, c0_n43_w116, c0_n43_w117, c0_n43_w118, c0_n43_w119, c0_n43_w120, c0_n43_w121, c0_n43_w122, c0_n43_w123, c0_n43_w124, c0_n43_w125, c0_n43_w126, c0_n43_w127, c0_n43_w128, c0_n43_w129, c0_n43_w130, c0_n43_w131, c0_n43_w132, c0_n43_w133, c0_n43_w134, c0_n43_w135, c0_n43_w136, c0_n43_w137, c0_n43_w138, c0_n43_w139, c0_n43_w140, c0_n43_w141, c0_n43_w142, c0_n43_w143, c0_n43_w144, c0_n43_w145, c0_n43_w146, c0_n43_w147, c0_n43_w148, c0_n43_w149, c0_n43_w150, c0_n43_w151, c0_n43_w152, c0_n43_w153, c0_n43_w154, c0_n43_w155, c0_n43_w156, c0_n43_w157, c0_n43_w158, c0_n43_w159, c0_n43_w160, c0_n43_w161, c0_n43_w162, c0_n43_w163, c0_n43_w164, c0_n43_w165, c0_n43_w166, c0_n43_w167, c0_n43_w168, c0_n43_w169, c0_n43_w170, c0_n43_w171, c0_n43_w172, c0_n43_w173, c0_n43_w174, c0_n43_w175, c0_n43_w176, c0_n43_w177, c0_n43_w178, c0_n43_w179, c0_n43_w180, c0_n43_w181, c0_n43_w182, c0_n43_w183, c0_n43_w184, c0_n43_w185, c0_n43_w186, c0_n43_w187, c0_n43_w188, c0_n43_w189, c0_n43_w190, c0_n43_w191, c0_n43_w192, c0_n43_w193, c0_n43_w194, c0_n43_w195, c0_n43_w196, c0_n43_w197, c0_n43_w198, c0_n43_w199, c0_n43_w200, c0_n44_w1, c0_n44_w2, c0_n44_w3, c0_n44_w4, c0_n44_w5, c0_n44_w6, c0_n44_w7, c0_n44_w8, c0_n44_w9, c0_n44_w10, c0_n44_w11, c0_n44_w12, c0_n44_w13, c0_n44_w14, c0_n44_w15, c0_n44_w16, c0_n44_w17, c0_n44_w18, c0_n44_w19, c0_n44_w20, c0_n44_w21, c0_n44_w22, c0_n44_w23, c0_n44_w24, c0_n44_w25, c0_n44_w26, c0_n44_w27, c0_n44_w28, c0_n44_w29, c0_n44_w30, c0_n44_w31, c0_n44_w32, c0_n44_w33, c0_n44_w34, c0_n44_w35, c0_n44_w36, c0_n44_w37, c0_n44_w38, c0_n44_w39, c0_n44_w40, c0_n44_w41, c0_n44_w42, c0_n44_w43, c0_n44_w44, c0_n44_w45, c0_n44_w46, c0_n44_w47, c0_n44_w48, c0_n44_w49, c0_n44_w50, c0_n44_w51, c0_n44_w52, c0_n44_w53, c0_n44_w54, c0_n44_w55, c0_n44_w56, c0_n44_w57, c0_n44_w58, c0_n44_w59, c0_n44_w60, c0_n44_w61, c0_n44_w62, c0_n44_w63, c0_n44_w64, c0_n44_w65, c0_n44_w66, c0_n44_w67, c0_n44_w68, c0_n44_w69, c0_n44_w70, c0_n44_w71, c0_n44_w72, c0_n44_w73, c0_n44_w74, c0_n44_w75, c0_n44_w76, c0_n44_w77, c0_n44_w78, c0_n44_w79, c0_n44_w80, c0_n44_w81, c0_n44_w82, c0_n44_w83, c0_n44_w84, c0_n44_w85, c0_n44_w86, c0_n44_w87, c0_n44_w88, c0_n44_w89, c0_n44_w90, c0_n44_w91, c0_n44_w92, c0_n44_w93, c0_n44_w94, c0_n44_w95, c0_n44_w96, c0_n44_w97, c0_n44_w98, c0_n44_w99, c0_n44_w100, c0_n44_w101, c0_n44_w102, c0_n44_w103, c0_n44_w104, c0_n44_w105, c0_n44_w106, c0_n44_w107, c0_n44_w108, c0_n44_w109, c0_n44_w110, c0_n44_w111, c0_n44_w112, c0_n44_w113, c0_n44_w114, c0_n44_w115, c0_n44_w116, c0_n44_w117, c0_n44_w118, c0_n44_w119, c0_n44_w120, c0_n44_w121, c0_n44_w122, c0_n44_w123, c0_n44_w124, c0_n44_w125, c0_n44_w126, c0_n44_w127, c0_n44_w128, c0_n44_w129, c0_n44_w130, c0_n44_w131, c0_n44_w132, c0_n44_w133, c0_n44_w134, c0_n44_w135, c0_n44_w136, c0_n44_w137, c0_n44_w138, c0_n44_w139, c0_n44_w140, c0_n44_w141, c0_n44_w142, c0_n44_w143, c0_n44_w144, c0_n44_w145, c0_n44_w146, c0_n44_w147, c0_n44_w148, c0_n44_w149, c0_n44_w150, c0_n44_w151, c0_n44_w152, c0_n44_w153, c0_n44_w154, c0_n44_w155, c0_n44_w156, c0_n44_w157, c0_n44_w158, c0_n44_w159, c0_n44_w160, c0_n44_w161, c0_n44_w162, c0_n44_w163, c0_n44_w164, c0_n44_w165, c0_n44_w166, c0_n44_w167, c0_n44_w168, c0_n44_w169, c0_n44_w170, c0_n44_w171, c0_n44_w172, c0_n44_w173, c0_n44_w174, c0_n44_w175, c0_n44_w176, c0_n44_w177, c0_n44_w178, c0_n44_w179, c0_n44_w180, c0_n44_w181, c0_n44_w182, c0_n44_w183, c0_n44_w184, c0_n44_w185, c0_n44_w186, c0_n44_w187, c0_n44_w188, c0_n44_w189, c0_n44_w190, c0_n44_w191, c0_n44_w192, c0_n44_w193, c0_n44_w194, c0_n44_w195, c0_n44_w196, c0_n44_w197, c0_n44_w198, c0_n44_w199, c0_n44_w200, c0_n45_w1, c0_n45_w2, c0_n45_w3, c0_n45_w4, c0_n45_w5, c0_n45_w6, c0_n45_w7, c0_n45_w8, c0_n45_w9, c0_n45_w10, c0_n45_w11, c0_n45_w12, c0_n45_w13, c0_n45_w14, c0_n45_w15, c0_n45_w16, c0_n45_w17, c0_n45_w18, c0_n45_w19, c0_n45_w20, c0_n45_w21, c0_n45_w22, c0_n45_w23, c0_n45_w24, c0_n45_w25, c0_n45_w26, c0_n45_w27, c0_n45_w28, c0_n45_w29, c0_n45_w30, c0_n45_w31, c0_n45_w32, c0_n45_w33, c0_n45_w34, c0_n45_w35, c0_n45_w36, c0_n45_w37, c0_n45_w38, c0_n45_w39, c0_n45_w40, c0_n45_w41, c0_n45_w42, c0_n45_w43, c0_n45_w44, c0_n45_w45, c0_n45_w46, c0_n45_w47, c0_n45_w48, c0_n45_w49, c0_n45_w50, c0_n45_w51, c0_n45_w52, c0_n45_w53, c0_n45_w54, c0_n45_w55, c0_n45_w56, c0_n45_w57, c0_n45_w58, c0_n45_w59, c0_n45_w60, c0_n45_w61, c0_n45_w62, c0_n45_w63, c0_n45_w64, c0_n45_w65, c0_n45_w66, c0_n45_w67, c0_n45_w68, c0_n45_w69, c0_n45_w70, c0_n45_w71, c0_n45_w72, c0_n45_w73, c0_n45_w74, c0_n45_w75, c0_n45_w76, c0_n45_w77, c0_n45_w78, c0_n45_w79, c0_n45_w80, c0_n45_w81, c0_n45_w82, c0_n45_w83, c0_n45_w84, c0_n45_w85, c0_n45_w86, c0_n45_w87, c0_n45_w88, c0_n45_w89, c0_n45_w90, c0_n45_w91, c0_n45_w92, c0_n45_w93, c0_n45_w94, c0_n45_w95, c0_n45_w96, c0_n45_w97, c0_n45_w98, c0_n45_w99, c0_n45_w100, c0_n45_w101, c0_n45_w102, c0_n45_w103, c0_n45_w104, c0_n45_w105, c0_n45_w106, c0_n45_w107, c0_n45_w108, c0_n45_w109, c0_n45_w110, c0_n45_w111, c0_n45_w112, c0_n45_w113, c0_n45_w114, c0_n45_w115, c0_n45_w116, c0_n45_w117, c0_n45_w118, c0_n45_w119, c0_n45_w120, c0_n45_w121, c0_n45_w122, c0_n45_w123, c0_n45_w124, c0_n45_w125, c0_n45_w126, c0_n45_w127, c0_n45_w128, c0_n45_w129, c0_n45_w130, c0_n45_w131, c0_n45_w132, c0_n45_w133, c0_n45_w134, c0_n45_w135, c0_n45_w136, c0_n45_w137, c0_n45_w138, c0_n45_w139, c0_n45_w140, c0_n45_w141, c0_n45_w142, c0_n45_w143, c0_n45_w144, c0_n45_w145, c0_n45_w146, c0_n45_w147, c0_n45_w148, c0_n45_w149, c0_n45_w150, c0_n45_w151, c0_n45_w152, c0_n45_w153, c0_n45_w154, c0_n45_w155, c0_n45_w156, c0_n45_w157, c0_n45_w158, c0_n45_w159, c0_n45_w160, c0_n45_w161, c0_n45_w162, c0_n45_w163, c0_n45_w164, c0_n45_w165, c0_n45_w166, c0_n45_w167, c0_n45_w168, c0_n45_w169, c0_n45_w170, c0_n45_w171, c0_n45_w172, c0_n45_w173, c0_n45_w174, c0_n45_w175, c0_n45_w176, c0_n45_w177, c0_n45_w178, c0_n45_w179, c0_n45_w180, c0_n45_w181, c0_n45_w182, c0_n45_w183, c0_n45_w184, c0_n45_w185, c0_n45_w186, c0_n45_w187, c0_n45_w188, c0_n45_w189, c0_n45_w190, c0_n45_w191, c0_n45_w192, c0_n45_w193, c0_n45_w194, c0_n45_w195, c0_n45_w196, c0_n45_w197, c0_n45_w198, c0_n45_w199, c0_n45_w200, c0_n46_w1, c0_n46_w2, c0_n46_w3, c0_n46_w4, c0_n46_w5, c0_n46_w6, c0_n46_w7, c0_n46_w8, c0_n46_w9, c0_n46_w10, c0_n46_w11, c0_n46_w12, c0_n46_w13, c0_n46_w14, c0_n46_w15, c0_n46_w16, c0_n46_w17, c0_n46_w18, c0_n46_w19, c0_n46_w20, c0_n46_w21, c0_n46_w22, c0_n46_w23, c0_n46_w24, c0_n46_w25, c0_n46_w26, c0_n46_w27, c0_n46_w28, c0_n46_w29, c0_n46_w30, c0_n46_w31, c0_n46_w32, c0_n46_w33, c0_n46_w34, c0_n46_w35, c0_n46_w36, c0_n46_w37, c0_n46_w38, c0_n46_w39, c0_n46_w40, c0_n46_w41, c0_n46_w42, c0_n46_w43, c0_n46_w44, c0_n46_w45, c0_n46_w46, c0_n46_w47, c0_n46_w48, c0_n46_w49, c0_n46_w50, c0_n46_w51, c0_n46_w52, c0_n46_w53, c0_n46_w54, c0_n46_w55, c0_n46_w56, c0_n46_w57, c0_n46_w58, c0_n46_w59, c0_n46_w60, c0_n46_w61, c0_n46_w62, c0_n46_w63, c0_n46_w64, c0_n46_w65, c0_n46_w66, c0_n46_w67, c0_n46_w68, c0_n46_w69, c0_n46_w70, c0_n46_w71, c0_n46_w72, c0_n46_w73, c0_n46_w74, c0_n46_w75, c0_n46_w76, c0_n46_w77, c0_n46_w78, c0_n46_w79, c0_n46_w80, c0_n46_w81, c0_n46_w82, c0_n46_w83, c0_n46_w84, c0_n46_w85, c0_n46_w86, c0_n46_w87, c0_n46_w88, c0_n46_w89, c0_n46_w90, c0_n46_w91, c0_n46_w92, c0_n46_w93, c0_n46_w94, c0_n46_w95, c0_n46_w96, c0_n46_w97, c0_n46_w98, c0_n46_w99, c0_n46_w100, c0_n46_w101, c0_n46_w102, c0_n46_w103, c0_n46_w104, c0_n46_w105, c0_n46_w106, c0_n46_w107, c0_n46_w108, c0_n46_w109, c0_n46_w110, c0_n46_w111, c0_n46_w112, c0_n46_w113, c0_n46_w114, c0_n46_w115, c0_n46_w116, c0_n46_w117, c0_n46_w118, c0_n46_w119, c0_n46_w120, c0_n46_w121, c0_n46_w122, c0_n46_w123, c0_n46_w124, c0_n46_w125, c0_n46_w126, c0_n46_w127, c0_n46_w128, c0_n46_w129, c0_n46_w130, c0_n46_w131, c0_n46_w132, c0_n46_w133, c0_n46_w134, c0_n46_w135, c0_n46_w136, c0_n46_w137, c0_n46_w138, c0_n46_w139, c0_n46_w140, c0_n46_w141, c0_n46_w142, c0_n46_w143, c0_n46_w144, c0_n46_w145, c0_n46_w146, c0_n46_w147, c0_n46_w148, c0_n46_w149, c0_n46_w150, c0_n46_w151, c0_n46_w152, c0_n46_w153, c0_n46_w154, c0_n46_w155, c0_n46_w156, c0_n46_w157, c0_n46_w158, c0_n46_w159, c0_n46_w160, c0_n46_w161, c0_n46_w162, c0_n46_w163, c0_n46_w164, c0_n46_w165, c0_n46_w166, c0_n46_w167, c0_n46_w168, c0_n46_w169, c0_n46_w170, c0_n46_w171, c0_n46_w172, c0_n46_w173, c0_n46_w174, c0_n46_w175, c0_n46_w176, c0_n46_w177, c0_n46_w178, c0_n46_w179, c0_n46_w180, c0_n46_w181, c0_n46_w182, c0_n46_w183, c0_n46_w184, c0_n46_w185, c0_n46_w186, c0_n46_w187, c0_n46_w188, c0_n46_w189, c0_n46_w190, c0_n46_w191, c0_n46_w192, c0_n46_w193, c0_n46_w194, c0_n46_w195, c0_n46_w196, c0_n46_w197, c0_n46_w198, c0_n46_w199, c0_n46_w200, c0_n47_w1, c0_n47_w2, c0_n47_w3, c0_n47_w4, c0_n47_w5, c0_n47_w6, c0_n47_w7, c0_n47_w8, c0_n47_w9, c0_n47_w10, c0_n47_w11, c0_n47_w12, c0_n47_w13, c0_n47_w14, c0_n47_w15, c0_n47_w16, c0_n47_w17, c0_n47_w18, c0_n47_w19, c0_n47_w20, c0_n47_w21, c0_n47_w22, c0_n47_w23, c0_n47_w24, c0_n47_w25, c0_n47_w26, c0_n47_w27, c0_n47_w28, c0_n47_w29, c0_n47_w30, c0_n47_w31, c0_n47_w32, c0_n47_w33, c0_n47_w34, c0_n47_w35, c0_n47_w36, c0_n47_w37, c0_n47_w38, c0_n47_w39, c0_n47_w40, c0_n47_w41, c0_n47_w42, c0_n47_w43, c0_n47_w44, c0_n47_w45, c0_n47_w46, c0_n47_w47, c0_n47_w48, c0_n47_w49, c0_n47_w50, c0_n47_w51, c0_n47_w52, c0_n47_w53, c0_n47_w54, c0_n47_w55, c0_n47_w56, c0_n47_w57, c0_n47_w58, c0_n47_w59, c0_n47_w60, c0_n47_w61, c0_n47_w62, c0_n47_w63, c0_n47_w64, c0_n47_w65, c0_n47_w66, c0_n47_w67, c0_n47_w68, c0_n47_w69, c0_n47_w70, c0_n47_w71, c0_n47_w72, c0_n47_w73, c0_n47_w74, c0_n47_w75, c0_n47_w76, c0_n47_w77, c0_n47_w78, c0_n47_w79, c0_n47_w80, c0_n47_w81, c0_n47_w82, c0_n47_w83, c0_n47_w84, c0_n47_w85, c0_n47_w86, c0_n47_w87, c0_n47_w88, c0_n47_w89, c0_n47_w90, c0_n47_w91, c0_n47_w92, c0_n47_w93, c0_n47_w94, c0_n47_w95, c0_n47_w96, c0_n47_w97, c0_n47_w98, c0_n47_w99, c0_n47_w100, c0_n47_w101, c0_n47_w102, c0_n47_w103, c0_n47_w104, c0_n47_w105, c0_n47_w106, c0_n47_w107, c0_n47_w108, c0_n47_w109, c0_n47_w110, c0_n47_w111, c0_n47_w112, c0_n47_w113, c0_n47_w114, c0_n47_w115, c0_n47_w116, c0_n47_w117, c0_n47_w118, c0_n47_w119, c0_n47_w120, c0_n47_w121, c0_n47_w122, c0_n47_w123, c0_n47_w124, c0_n47_w125, c0_n47_w126, c0_n47_w127, c0_n47_w128, c0_n47_w129, c0_n47_w130, c0_n47_w131, c0_n47_w132, c0_n47_w133, c0_n47_w134, c0_n47_w135, c0_n47_w136, c0_n47_w137, c0_n47_w138, c0_n47_w139, c0_n47_w140, c0_n47_w141, c0_n47_w142, c0_n47_w143, c0_n47_w144, c0_n47_w145, c0_n47_w146, c0_n47_w147, c0_n47_w148, c0_n47_w149, c0_n47_w150, c0_n47_w151, c0_n47_w152, c0_n47_w153, c0_n47_w154, c0_n47_w155, c0_n47_w156, c0_n47_w157, c0_n47_w158, c0_n47_w159, c0_n47_w160, c0_n47_w161, c0_n47_w162, c0_n47_w163, c0_n47_w164, c0_n47_w165, c0_n47_w166, c0_n47_w167, c0_n47_w168, c0_n47_w169, c0_n47_w170, c0_n47_w171, c0_n47_w172, c0_n47_w173, c0_n47_w174, c0_n47_w175, c0_n47_w176, c0_n47_w177, c0_n47_w178, c0_n47_w179, c0_n47_w180, c0_n47_w181, c0_n47_w182, c0_n47_w183, c0_n47_w184, c0_n47_w185, c0_n47_w186, c0_n47_w187, c0_n47_w188, c0_n47_w189, c0_n47_w190, c0_n47_w191, c0_n47_w192, c0_n47_w193, c0_n47_w194, c0_n47_w195, c0_n47_w196, c0_n47_w197, c0_n47_w198, c0_n47_w199, c0_n47_w200, c0_n48_w1, c0_n48_w2, c0_n48_w3, c0_n48_w4, c0_n48_w5, c0_n48_w6, c0_n48_w7, c0_n48_w8, c0_n48_w9, c0_n48_w10, c0_n48_w11, c0_n48_w12, c0_n48_w13, c0_n48_w14, c0_n48_w15, c0_n48_w16, c0_n48_w17, c0_n48_w18, c0_n48_w19, c0_n48_w20, c0_n48_w21, c0_n48_w22, c0_n48_w23, c0_n48_w24, c0_n48_w25, c0_n48_w26, c0_n48_w27, c0_n48_w28, c0_n48_w29, c0_n48_w30, c0_n48_w31, c0_n48_w32, c0_n48_w33, c0_n48_w34, c0_n48_w35, c0_n48_w36, c0_n48_w37, c0_n48_w38, c0_n48_w39, c0_n48_w40, c0_n48_w41, c0_n48_w42, c0_n48_w43, c0_n48_w44, c0_n48_w45, c0_n48_w46, c0_n48_w47, c0_n48_w48, c0_n48_w49, c0_n48_w50, c0_n48_w51, c0_n48_w52, c0_n48_w53, c0_n48_w54, c0_n48_w55, c0_n48_w56, c0_n48_w57, c0_n48_w58, c0_n48_w59, c0_n48_w60, c0_n48_w61, c0_n48_w62, c0_n48_w63, c0_n48_w64, c0_n48_w65, c0_n48_w66, c0_n48_w67, c0_n48_w68, c0_n48_w69, c0_n48_w70, c0_n48_w71, c0_n48_w72, c0_n48_w73, c0_n48_w74, c0_n48_w75, c0_n48_w76, c0_n48_w77, c0_n48_w78, c0_n48_w79, c0_n48_w80, c0_n48_w81, c0_n48_w82, c0_n48_w83, c0_n48_w84, c0_n48_w85, c0_n48_w86, c0_n48_w87, c0_n48_w88, c0_n48_w89, c0_n48_w90, c0_n48_w91, c0_n48_w92, c0_n48_w93, c0_n48_w94, c0_n48_w95, c0_n48_w96, c0_n48_w97, c0_n48_w98, c0_n48_w99, c0_n48_w100, c0_n48_w101, c0_n48_w102, c0_n48_w103, c0_n48_w104, c0_n48_w105, c0_n48_w106, c0_n48_w107, c0_n48_w108, c0_n48_w109, c0_n48_w110, c0_n48_w111, c0_n48_w112, c0_n48_w113, c0_n48_w114, c0_n48_w115, c0_n48_w116, c0_n48_w117, c0_n48_w118, c0_n48_w119, c0_n48_w120, c0_n48_w121, c0_n48_w122, c0_n48_w123, c0_n48_w124, c0_n48_w125, c0_n48_w126, c0_n48_w127, c0_n48_w128, c0_n48_w129, c0_n48_w130, c0_n48_w131, c0_n48_w132, c0_n48_w133, c0_n48_w134, c0_n48_w135, c0_n48_w136, c0_n48_w137, c0_n48_w138, c0_n48_w139, c0_n48_w140, c0_n48_w141, c0_n48_w142, c0_n48_w143, c0_n48_w144, c0_n48_w145, c0_n48_w146, c0_n48_w147, c0_n48_w148, c0_n48_w149, c0_n48_w150, c0_n48_w151, c0_n48_w152, c0_n48_w153, c0_n48_w154, c0_n48_w155, c0_n48_w156, c0_n48_w157, c0_n48_w158, c0_n48_w159, c0_n48_w160, c0_n48_w161, c0_n48_w162, c0_n48_w163, c0_n48_w164, c0_n48_w165, c0_n48_w166, c0_n48_w167, c0_n48_w168, c0_n48_w169, c0_n48_w170, c0_n48_w171, c0_n48_w172, c0_n48_w173, c0_n48_w174, c0_n48_w175, c0_n48_w176, c0_n48_w177, c0_n48_w178, c0_n48_w179, c0_n48_w180, c0_n48_w181, c0_n48_w182, c0_n48_w183, c0_n48_w184, c0_n48_w185, c0_n48_w186, c0_n48_w187, c0_n48_w188, c0_n48_w189, c0_n48_w190, c0_n48_w191, c0_n48_w192, c0_n48_w193, c0_n48_w194, c0_n48_w195, c0_n48_w196, c0_n48_w197, c0_n48_w198, c0_n48_w199, c0_n48_w200, c0_n49_w1, c0_n49_w2, c0_n49_w3, c0_n49_w4, c0_n49_w5, c0_n49_w6, c0_n49_w7, c0_n49_w8, c0_n49_w9, c0_n49_w10, c0_n49_w11, c0_n49_w12, c0_n49_w13, c0_n49_w14, c0_n49_w15, c0_n49_w16, c0_n49_w17, c0_n49_w18, c0_n49_w19, c0_n49_w20, c0_n49_w21, c0_n49_w22, c0_n49_w23, c0_n49_w24, c0_n49_w25, c0_n49_w26, c0_n49_w27, c0_n49_w28, c0_n49_w29, c0_n49_w30, c0_n49_w31, c0_n49_w32, c0_n49_w33, c0_n49_w34, c0_n49_w35, c0_n49_w36, c0_n49_w37, c0_n49_w38, c0_n49_w39, c0_n49_w40, c0_n49_w41, c0_n49_w42, c0_n49_w43, c0_n49_w44, c0_n49_w45, c0_n49_w46, c0_n49_w47, c0_n49_w48, c0_n49_w49, c0_n49_w50, c0_n49_w51, c0_n49_w52, c0_n49_w53, c0_n49_w54, c0_n49_w55, c0_n49_w56, c0_n49_w57, c0_n49_w58, c0_n49_w59, c0_n49_w60, c0_n49_w61, c0_n49_w62, c0_n49_w63, c0_n49_w64, c0_n49_w65, c0_n49_w66, c0_n49_w67, c0_n49_w68, c0_n49_w69, c0_n49_w70, c0_n49_w71, c0_n49_w72, c0_n49_w73, c0_n49_w74, c0_n49_w75, c0_n49_w76, c0_n49_w77, c0_n49_w78, c0_n49_w79, c0_n49_w80, c0_n49_w81, c0_n49_w82, c0_n49_w83, c0_n49_w84, c0_n49_w85, c0_n49_w86, c0_n49_w87, c0_n49_w88, c0_n49_w89, c0_n49_w90, c0_n49_w91, c0_n49_w92, c0_n49_w93, c0_n49_w94, c0_n49_w95, c0_n49_w96, c0_n49_w97, c0_n49_w98, c0_n49_w99, c0_n49_w100, c0_n49_w101, c0_n49_w102, c0_n49_w103, c0_n49_w104, c0_n49_w105, c0_n49_w106, c0_n49_w107, c0_n49_w108, c0_n49_w109, c0_n49_w110, c0_n49_w111, c0_n49_w112, c0_n49_w113, c0_n49_w114, c0_n49_w115, c0_n49_w116, c0_n49_w117, c0_n49_w118, c0_n49_w119, c0_n49_w120, c0_n49_w121, c0_n49_w122, c0_n49_w123, c0_n49_w124, c0_n49_w125, c0_n49_w126, c0_n49_w127, c0_n49_w128, c0_n49_w129, c0_n49_w130, c0_n49_w131, c0_n49_w132, c0_n49_w133, c0_n49_w134, c0_n49_w135, c0_n49_w136, c0_n49_w137, c0_n49_w138, c0_n49_w139, c0_n49_w140, c0_n49_w141, c0_n49_w142, c0_n49_w143, c0_n49_w144, c0_n49_w145, c0_n49_w146, c0_n49_w147, c0_n49_w148, c0_n49_w149, c0_n49_w150, c0_n49_w151, c0_n49_w152, c0_n49_w153, c0_n49_w154, c0_n49_w155, c0_n49_w156, c0_n49_w157, c0_n49_w158, c0_n49_w159, c0_n49_w160, c0_n49_w161, c0_n49_w162, c0_n49_w163, c0_n49_w164, c0_n49_w165, c0_n49_w166, c0_n49_w167, c0_n49_w168, c0_n49_w169, c0_n49_w170, c0_n49_w171, c0_n49_w172, c0_n49_w173, c0_n49_w174, c0_n49_w175, c0_n49_w176, c0_n49_w177, c0_n49_w178, c0_n49_w179, c0_n49_w180, c0_n49_w181, c0_n49_w182, c0_n49_w183, c0_n49_w184, c0_n49_w185, c0_n49_w186, c0_n49_w187, c0_n49_w188, c0_n49_w189, c0_n49_w190, c0_n49_w191, c0_n49_w192, c0_n49_w193, c0_n49_w194, c0_n49_w195, c0_n49_w196, c0_n49_w197, c0_n49_w198, c0_n49_w199, c0_n49_w200, c0_n50_w1, c0_n50_w2, c0_n50_w3, c0_n50_w4, c0_n50_w5, c0_n50_w6, c0_n50_w7, c0_n50_w8, c0_n50_w9, c0_n50_w10, c0_n50_w11, c0_n50_w12, c0_n50_w13, c0_n50_w14, c0_n50_w15, c0_n50_w16, c0_n50_w17, c0_n50_w18, c0_n50_w19, c0_n50_w20, c0_n50_w21, c0_n50_w22, c0_n50_w23, c0_n50_w24, c0_n50_w25, c0_n50_w26, c0_n50_w27, c0_n50_w28, c0_n50_w29, c0_n50_w30, c0_n50_w31, c0_n50_w32, c0_n50_w33, c0_n50_w34, c0_n50_w35, c0_n50_w36, c0_n50_w37, c0_n50_w38, c0_n50_w39, c0_n50_w40, c0_n50_w41, c0_n50_w42, c0_n50_w43, c0_n50_w44, c0_n50_w45, c0_n50_w46, c0_n50_w47, c0_n50_w48, c0_n50_w49, c0_n50_w50, c0_n50_w51, c0_n50_w52, c0_n50_w53, c0_n50_w54, c0_n50_w55, c0_n50_w56, c0_n50_w57, c0_n50_w58, c0_n50_w59, c0_n50_w60, c0_n50_w61, c0_n50_w62, c0_n50_w63, c0_n50_w64, c0_n50_w65, c0_n50_w66, c0_n50_w67, c0_n50_w68, c0_n50_w69, c0_n50_w70, c0_n50_w71, c0_n50_w72, c0_n50_w73, c0_n50_w74, c0_n50_w75, c0_n50_w76, c0_n50_w77, c0_n50_w78, c0_n50_w79, c0_n50_w80, c0_n50_w81, c0_n50_w82, c0_n50_w83, c0_n50_w84, c0_n50_w85, c0_n50_w86, c0_n50_w87, c0_n50_w88, c0_n50_w89, c0_n50_w90, c0_n50_w91, c0_n50_w92, c0_n50_w93, c0_n50_w94, c0_n50_w95, c0_n50_w96, c0_n50_w97, c0_n50_w98, c0_n50_w99, c0_n50_w100, c0_n50_w101, c0_n50_w102, c0_n50_w103, c0_n50_w104, c0_n50_w105, c0_n50_w106, c0_n50_w107, c0_n50_w108, c0_n50_w109, c0_n50_w110, c0_n50_w111, c0_n50_w112, c0_n50_w113, c0_n50_w114, c0_n50_w115, c0_n50_w116, c0_n50_w117, c0_n50_w118, c0_n50_w119, c0_n50_w120, c0_n50_w121, c0_n50_w122, c0_n50_w123, c0_n50_w124, c0_n50_w125, c0_n50_w126, c0_n50_w127, c0_n50_w128, c0_n50_w129, c0_n50_w130, c0_n50_w131, c0_n50_w132, c0_n50_w133, c0_n50_w134, c0_n50_w135, c0_n50_w136, c0_n50_w137, c0_n50_w138, c0_n50_w139, c0_n50_w140, c0_n50_w141, c0_n50_w142, c0_n50_w143, c0_n50_w144, c0_n50_w145, c0_n50_w146, c0_n50_w147, c0_n50_w148, c0_n50_w149, c0_n50_w150, c0_n50_w151, c0_n50_w152, c0_n50_w153, c0_n50_w154, c0_n50_w155, c0_n50_w156, c0_n50_w157, c0_n50_w158, c0_n50_w159, c0_n50_w160, c0_n50_w161, c0_n50_w162, c0_n50_w163, c0_n50_w164, c0_n50_w165, c0_n50_w166, c0_n50_w167, c0_n50_w168, c0_n50_w169, c0_n50_w170, c0_n50_w171, c0_n50_w172, c0_n50_w173, c0_n50_w174, c0_n50_w175, c0_n50_w176, c0_n50_w177, c0_n50_w178, c0_n50_w179, c0_n50_w180, c0_n50_w181, c0_n50_w182, c0_n50_w183, c0_n50_w184, c0_n50_w185, c0_n50_w186, c0_n50_w187, c0_n50_w188, c0_n50_w189, c0_n50_w190, c0_n50_w191, c0_n50_w192, c0_n50_w193, c0_n50_w194, c0_n50_w195, c0_n50_w196, c0_n50_w197, c0_n50_w198, c0_n50_w199, c0_n50_w200, c0_n51_w1, c0_n51_w2, c0_n51_w3, c0_n51_w4, c0_n51_w5, c0_n51_w6, c0_n51_w7, c0_n51_w8, c0_n51_w9, c0_n51_w10, c0_n51_w11, c0_n51_w12, c0_n51_w13, c0_n51_w14, c0_n51_w15, c0_n51_w16, c0_n51_w17, c0_n51_w18, c0_n51_w19, c0_n51_w20, c0_n51_w21, c0_n51_w22, c0_n51_w23, c0_n51_w24, c0_n51_w25, c0_n51_w26, c0_n51_w27, c0_n51_w28, c0_n51_w29, c0_n51_w30, c0_n51_w31, c0_n51_w32, c0_n51_w33, c0_n51_w34, c0_n51_w35, c0_n51_w36, c0_n51_w37, c0_n51_w38, c0_n51_w39, c0_n51_w40, c0_n51_w41, c0_n51_w42, c0_n51_w43, c0_n51_w44, c0_n51_w45, c0_n51_w46, c0_n51_w47, c0_n51_w48, c0_n51_w49, c0_n51_w50, c0_n51_w51, c0_n51_w52, c0_n51_w53, c0_n51_w54, c0_n51_w55, c0_n51_w56, c0_n51_w57, c0_n51_w58, c0_n51_w59, c0_n51_w60, c0_n51_w61, c0_n51_w62, c0_n51_w63, c0_n51_w64, c0_n51_w65, c0_n51_w66, c0_n51_w67, c0_n51_w68, c0_n51_w69, c0_n51_w70, c0_n51_w71, c0_n51_w72, c0_n51_w73, c0_n51_w74, c0_n51_w75, c0_n51_w76, c0_n51_w77, c0_n51_w78, c0_n51_w79, c0_n51_w80, c0_n51_w81, c0_n51_w82, c0_n51_w83, c0_n51_w84, c0_n51_w85, c0_n51_w86, c0_n51_w87, c0_n51_w88, c0_n51_w89, c0_n51_w90, c0_n51_w91, c0_n51_w92, c0_n51_w93, c0_n51_w94, c0_n51_w95, c0_n51_w96, c0_n51_w97, c0_n51_w98, c0_n51_w99, c0_n51_w100, c0_n51_w101, c0_n51_w102, c0_n51_w103, c0_n51_w104, c0_n51_w105, c0_n51_w106, c0_n51_w107, c0_n51_w108, c0_n51_w109, c0_n51_w110, c0_n51_w111, c0_n51_w112, c0_n51_w113, c0_n51_w114, c0_n51_w115, c0_n51_w116, c0_n51_w117, c0_n51_w118, c0_n51_w119, c0_n51_w120, c0_n51_w121, c0_n51_w122, c0_n51_w123, c0_n51_w124, c0_n51_w125, c0_n51_w126, c0_n51_w127, c0_n51_w128, c0_n51_w129, c0_n51_w130, c0_n51_w131, c0_n51_w132, c0_n51_w133, c0_n51_w134, c0_n51_w135, c0_n51_w136, c0_n51_w137, c0_n51_w138, c0_n51_w139, c0_n51_w140, c0_n51_w141, c0_n51_w142, c0_n51_w143, c0_n51_w144, c0_n51_w145, c0_n51_w146, c0_n51_w147, c0_n51_w148, c0_n51_w149, c0_n51_w150, c0_n51_w151, c0_n51_w152, c0_n51_w153, c0_n51_w154, c0_n51_w155, c0_n51_w156, c0_n51_w157, c0_n51_w158, c0_n51_w159, c0_n51_w160, c0_n51_w161, c0_n51_w162, c0_n51_w163, c0_n51_w164, c0_n51_w165, c0_n51_w166, c0_n51_w167, c0_n51_w168, c0_n51_w169, c0_n51_w170, c0_n51_w171, c0_n51_w172, c0_n51_w173, c0_n51_w174, c0_n51_w175, c0_n51_w176, c0_n51_w177, c0_n51_w178, c0_n51_w179, c0_n51_w180, c0_n51_w181, c0_n51_w182, c0_n51_w183, c0_n51_w184, c0_n51_w185, c0_n51_w186, c0_n51_w187, c0_n51_w188, c0_n51_w189, c0_n51_w190, c0_n51_w191, c0_n51_w192, c0_n51_w193, c0_n51_w194, c0_n51_w195, c0_n51_w196, c0_n51_w197, c0_n51_w198, c0_n51_w199, c0_n51_w200, c0_n52_w1, c0_n52_w2, c0_n52_w3, c0_n52_w4, c0_n52_w5, c0_n52_w6, c0_n52_w7, c0_n52_w8, c0_n52_w9, c0_n52_w10, c0_n52_w11, c0_n52_w12, c0_n52_w13, c0_n52_w14, c0_n52_w15, c0_n52_w16, c0_n52_w17, c0_n52_w18, c0_n52_w19, c0_n52_w20, c0_n52_w21, c0_n52_w22, c0_n52_w23, c0_n52_w24, c0_n52_w25, c0_n52_w26, c0_n52_w27, c0_n52_w28, c0_n52_w29, c0_n52_w30, c0_n52_w31, c0_n52_w32, c0_n52_w33, c0_n52_w34, c0_n52_w35, c0_n52_w36, c0_n52_w37, c0_n52_w38, c0_n52_w39, c0_n52_w40, c0_n52_w41, c0_n52_w42, c0_n52_w43, c0_n52_w44, c0_n52_w45, c0_n52_w46, c0_n52_w47, c0_n52_w48, c0_n52_w49, c0_n52_w50, c0_n52_w51, c0_n52_w52, c0_n52_w53, c0_n52_w54, c0_n52_w55, c0_n52_w56, c0_n52_w57, c0_n52_w58, c0_n52_w59, c0_n52_w60, c0_n52_w61, c0_n52_w62, c0_n52_w63, c0_n52_w64, c0_n52_w65, c0_n52_w66, c0_n52_w67, c0_n52_w68, c0_n52_w69, c0_n52_w70, c0_n52_w71, c0_n52_w72, c0_n52_w73, c0_n52_w74, c0_n52_w75, c0_n52_w76, c0_n52_w77, c0_n52_w78, c0_n52_w79, c0_n52_w80, c0_n52_w81, c0_n52_w82, c0_n52_w83, c0_n52_w84, c0_n52_w85, c0_n52_w86, c0_n52_w87, c0_n52_w88, c0_n52_w89, c0_n52_w90, c0_n52_w91, c0_n52_w92, c0_n52_w93, c0_n52_w94, c0_n52_w95, c0_n52_w96, c0_n52_w97, c0_n52_w98, c0_n52_w99, c0_n52_w100, c0_n52_w101, c0_n52_w102, c0_n52_w103, c0_n52_w104, c0_n52_w105, c0_n52_w106, c0_n52_w107, c0_n52_w108, c0_n52_w109, c0_n52_w110, c0_n52_w111, c0_n52_w112, c0_n52_w113, c0_n52_w114, c0_n52_w115, c0_n52_w116, c0_n52_w117, c0_n52_w118, c0_n52_w119, c0_n52_w120, c0_n52_w121, c0_n52_w122, c0_n52_w123, c0_n52_w124, c0_n52_w125, c0_n52_w126, c0_n52_w127, c0_n52_w128, c0_n52_w129, c0_n52_w130, c0_n52_w131, c0_n52_w132, c0_n52_w133, c0_n52_w134, c0_n52_w135, c0_n52_w136, c0_n52_w137, c0_n52_w138, c0_n52_w139, c0_n52_w140, c0_n52_w141, c0_n52_w142, c0_n52_w143, c0_n52_w144, c0_n52_w145, c0_n52_w146, c0_n52_w147, c0_n52_w148, c0_n52_w149, c0_n52_w150, c0_n52_w151, c0_n52_w152, c0_n52_w153, c0_n52_w154, c0_n52_w155, c0_n52_w156, c0_n52_w157, c0_n52_w158, c0_n52_w159, c0_n52_w160, c0_n52_w161, c0_n52_w162, c0_n52_w163, c0_n52_w164, c0_n52_w165, c0_n52_w166, c0_n52_w167, c0_n52_w168, c0_n52_w169, c0_n52_w170, c0_n52_w171, c0_n52_w172, c0_n52_w173, c0_n52_w174, c0_n52_w175, c0_n52_w176, c0_n52_w177, c0_n52_w178, c0_n52_w179, c0_n52_w180, c0_n52_w181, c0_n52_w182, c0_n52_w183, c0_n52_w184, c0_n52_w185, c0_n52_w186, c0_n52_w187, c0_n52_w188, c0_n52_w189, c0_n52_w190, c0_n52_w191, c0_n52_w192, c0_n52_w193, c0_n52_w194, c0_n52_w195, c0_n52_w196, c0_n52_w197, c0_n52_w198, c0_n52_w199, c0_n52_w200, c0_n53_w1, c0_n53_w2, c0_n53_w3, c0_n53_w4, c0_n53_w5, c0_n53_w6, c0_n53_w7, c0_n53_w8, c0_n53_w9, c0_n53_w10, c0_n53_w11, c0_n53_w12, c0_n53_w13, c0_n53_w14, c0_n53_w15, c0_n53_w16, c0_n53_w17, c0_n53_w18, c0_n53_w19, c0_n53_w20, c0_n53_w21, c0_n53_w22, c0_n53_w23, c0_n53_w24, c0_n53_w25, c0_n53_w26, c0_n53_w27, c0_n53_w28, c0_n53_w29, c0_n53_w30, c0_n53_w31, c0_n53_w32, c0_n53_w33, c0_n53_w34, c0_n53_w35, c0_n53_w36, c0_n53_w37, c0_n53_w38, c0_n53_w39, c0_n53_w40, c0_n53_w41, c0_n53_w42, c0_n53_w43, c0_n53_w44, c0_n53_w45, c0_n53_w46, c0_n53_w47, c0_n53_w48, c0_n53_w49, c0_n53_w50, c0_n53_w51, c0_n53_w52, c0_n53_w53, c0_n53_w54, c0_n53_w55, c0_n53_w56, c0_n53_w57, c0_n53_w58, c0_n53_w59, c0_n53_w60, c0_n53_w61, c0_n53_w62, c0_n53_w63, c0_n53_w64, c0_n53_w65, c0_n53_w66, c0_n53_w67, c0_n53_w68, c0_n53_w69, c0_n53_w70, c0_n53_w71, c0_n53_w72, c0_n53_w73, c0_n53_w74, c0_n53_w75, c0_n53_w76, c0_n53_w77, c0_n53_w78, c0_n53_w79, c0_n53_w80, c0_n53_w81, c0_n53_w82, c0_n53_w83, c0_n53_w84, c0_n53_w85, c0_n53_w86, c0_n53_w87, c0_n53_w88, c0_n53_w89, c0_n53_w90, c0_n53_w91, c0_n53_w92, c0_n53_w93, c0_n53_w94, c0_n53_w95, c0_n53_w96, c0_n53_w97, c0_n53_w98, c0_n53_w99, c0_n53_w100, c0_n53_w101, c0_n53_w102, c0_n53_w103, c0_n53_w104, c0_n53_w105, c0_n53_w106, c0_n53_w107, c0_n53_w108, c0_n53_w109, c0_n53_w110, c0_n53_w111, c0_n53_w112, c0_n53_w113, c0_n53_w114, c0_n53_w115, c0_n53_w116, c0_n53_w117, c0_n53_w118, c0_n53_w119, c0_n53_w120, c0_n53_w121, c0_n53_w122, c0_n53_w123, c0_n53_w124, c0_n53_w125, c0_n53_w126, c0_n53_w127, c0_n53_w128, c0_n53_w129, c0_n53_w130, c0_n53_w131, c0_n53_w132, c0_n53_w133, c0_n53_w134, c0_n53_w135, c0_n53_w136, c0_n53_w137, c0_n53_w138, c0_n53_w139, c0_n53_w140, c0_n53_w141, c0_n53_w142, c0_n53_w143, c0_n53_w144, c0_n53_w145, c0_n53_w146, c0_n53_w147, c0_n53_w148, c0_n53_w149, c0_n53_w150, c0_n53_w151, c0_n53_w152, c0_n53_w153, c0_n53_w154, c0_n53_w155, c0_n53_w156, c0_n53_w157, c0_n53_w158, c0_n53_w159, c0_n53_w160, c0_n53_w161, c0_n53_w162, c0_n53_w163, c0_n53_w164, c0_n53_w165, c0_n53_w166, c0_n53_w167, c0_n53_w168, c0_n53_w169, c0_n53_w170, c0_n53_w171, c0_n53_w172, c0_n53_w173, c0_n53_w174, c0_n53_w175, c0_n53_w176, c0_n53_w177, c0_n53_w178, c0_n53_w179, c0_n53_w180, c0_n53_w181, c0_n53_w182, c0_n53_w183, c0_n53_w184, c0_n53_w185, c0_n53_w186, c0_n53_w187, c0_n53_w188, c0_n53_w189, c0_n53_w190, c0_n53_w191, c0_n53_w192, c0_n53_w193, c0_n53_w194, c0_n53_w195, c0_n53_w196, c0_n53_w197, c0_n53_w198, c0_n53_w199, c0_n53_w200, c0_n54_w1, c0_n54_w2, c0_n54_w3, c0_n54_w4, c0_n54_w5, c0_n54_w6, c0_n54_w7, c0_n54_w8, c0_n54_w9, c0_n54_w10, c0_n54_w11, c0_n54_w12, c0_n54_w13, c0_n54_w14, c0_n54_w15, c0_n54_w16, c0_n54_w17, c0_n54_w18, c0_n54_w19, c0_n54_w20, c0_n54_w21, c0_n54_w22, c0_n54_w23, c0_n54_w24, c0_n54_w25, c0_n54_w26, c0_n54_w27, c0_n54_w28, c0_n54_w29, c0_n54_w30, c0_n54_w31, c0_n54_w32, c0_n54_w33, c0_n54_w34, c0_n54_w35, c0_n54_w36, c0_n54_w37, c0_n54_w38, c0_n54_w39, c0_n54_w40, c0_n54_w41, c0_n54_w42, c0_n54_w43, c0_n54_w44, c0_n54_w45, c0_n54_w46, c0_n54_w47, c0_n54_w48, c0_n54_w49, c0_n54_w50, c0_n54_w51, c0_n54_w52, c0_n54_w53, c0_n54_w54, c0_n54_w55, c0_n54_w56, c0_n54_w57, c0_n54_w58, c0_n54_w59, c0_n54_w60, c0_n54_w61, c0_n54_w62, c0_n54_w63, c0_n54_w64, c0_n54_w65, c0_n54_w66, c0_n54_w67, c0_n54_w68, c0_n54_w69, c0_n54_w70, c0_n54_w71, c0_n54_w72, c0_n54_w73, c0_n54_w74, c0_n54_w75, c0_n54_w76, c0_n54_w77, c0_n54_w78, c0_n54_w79, c0_n54_w80, c0_n54_w81, c0_n54_w82, c0_n54_w83, c0_n54_w84, c0_n54_w85, c0_n54_w86, c0_n54_w87, c0_n54_w88, c0_n54_w89, c0_n54_w90, c0_n54_w91, c0_n54_w92, c0_n54_w93, c0_n54_w94, c0_n54_w95, c0_n54_w96, c0_n54_w97, c0_n54_w98, c0_n54_w99, c0_n54_w100, c0_n54_w101, c0_n54_w102, c0_n54_w103, c0_n54_w104, c0_n54_w105, c0_n54_w106, c0_n54_w107, c0_n54_w108, c0_n54_w109, c0_n54_w110, c0_n54_w111, c0_n54_w112, c0_n54_w113, c0_n54_w114, c0_n54_w115, c0_n54_w116, c0_n54_w117, c0_n54_w118, c0_n54_w119, c0_n54_w120, c0_n54_w121, c0_n54_w122, c0_n54_w123, c0_n54_w124, c0_n54_w125, c0_n54_w126, c0_n54_w127, c0_n54_w128, c0_n54_w129, c0_n54_w130, c0_n54_w131, c0_n54_w132, c0_n54_w133, c0_n54_w134, c0_n54_w135, c0_n54_w136, c0_n54_w137, c0_n54_w138, c0_n54_w139, c0_n54_w140, c0_n54_w141, c0_n54_w142, c0_n54_w143, c0_n54_w144, c0_n54_w145, c0_n54_w146, c0_n54_w147, c0_n54_w148, c0_n54_w149, c0_n54_w150, c0_n54_w151, c0_n54_w152, c0_n54_w153, c0_n54_w154, c0_n54_w155, c0_n54_w156, c0_n54_w157, c0_n54_w158, c0_n54_w159, c0_n54_w160, c0_n54_w161, c0_n54_w162, c0_n54_w163, c0_n54_w164, c0_n54_w165, c0_n54_w166, c0_n54_w167, c0_n54_w168, c0_n54_w169, c0_n54_w170, c0_n54_w171, c0_n54_w172, c0_n54_w173, c0_n54_w174, c0_n54_w175, c0_n54_w176, c0_n54_w177, c0_n54_w178, c0_n54_w179, c0_n54_w180, c0_n54_w181, c0_n54_w182, c0_n54_w183, c0_n54_w184, c0_n54_w185, c0_n54_w186, c0_n54_w187, c0_n54_w188, c0_n54_w189, c0_n54_w190, c0_n54_w191, c0_n54_w192, c0_n54_w193, c0_n54_w194, c0_n54_w195, c0_n54_w196, c0_n54_w197, c0_n54_w198, c0_n54_w199, c0_n54_w200, c0_n55_w1, c0_n55_w2, c0_n55_w3, c0_n55_w4, c0_n55_w5, c0_n55_w6, c0_n55_w7, c0_n55_w8, c0_n55_w9, c0_n55_w10, c0_n55_w11, c0_n55_w12, c0_n55_w13, c0_n55_w14, c0_n55_w15, c0_n55_w16, c0_n55_w17, c0_n55_w18, c0_n55_w19, c0_n55_w20, c0_n55_w21, c0_n55_w22, c0_n55_w23, c0_n55_w24, c0_n55_w25, c0_n55_w26, c0_n55_w27, c0_n55_w28, c0_n55_w29, c0_n55_w30, c0_n55_w31, c0_n55_w32, c0_n55_w33, c0_n55_w34, c0_n55_w35, c0_n55_w36, c0_n55_w37, c0_n55_w38, c0_n55_w39, c0_n55_w40, c0_n55_w41, c0_n55_w42, c0_n55_w43, c0_n55_w44, c0_n55_w45, c0_n55_w46, c0_n55_w47, c0_n55_w48, c0_n55_w49, c0_n55_w50, c0_n55_w51, c0_n55_w52, c0_n55_w53, c0_n55_w54, c0_n55_w55, c0_n55_w56, c0_n55_w57, c0_n55_w58, c0_n55_w59, c0_n55_w60, c0_n55_w61, c0_n55_w62, c0_n55_w63, c0_n55_w64, c0_n55_w65, c0_n55_w66, c0_n55_w67, c0_n55_w68, c0_n55_w69, c0_n55_w70, c0_n55_w71, c0_n55_w72, c0_n55_w73, c0_n55_w74, c0_n55_w75, c0_n55_w76, c0_n55_w77, c0_n55_w78, c0_n55_w79, c0_n55_w80, c0_n55_w81, c0_n55_w82, c0_n55_w83, c0_n55_w84, c0_n55_w85, c0_n55_w86, c0_n55_w87, c0_n55_w88, c0_n55_w89, c0_n55_w90, c0_n55_w91, c0_n55_w92, c0_n55_w93, c0_n55_w94, c0_n55_w95, c0_n55_w96, c0_n55_w97, c0_n55_w98, c0_n55_w99, c0_n55_w100, c0_n55_w101, c0_n55_w102, c0_n55_w103, c0_n55_w104, c0_n55_w105, c0_n55_w106, c0_n55_w107, c0_n55_w108, c0_n55_w109, c0_n55_w110, c0_n55_w111, c0_n55_w112, c0_n55_w113, c0_n55_w114, c0_n55_w115, c0_n55_w116, c0_n55_w117, c0_n55_w118, c0_n55_w119, c0_n55_w120, c0_n55_w121, c0_n55_w122, c0_n55_w123, c0_n55_w124, c0_n55_w125, c0_n55_w126, c0_n55_w127, c0_n55_w128, c0_n55_w129, c0_n55_w130, c0_n55_w131, c0_n55_w132, c0_n55_w133, c0_n55_w134, c0_n55_w135, c0_n55_w136, c0_n55_w137, c0_n55_w138, c0_n55_w139, c0_n55_w140, c0_n55_w141, c0_n55_w142, c0_n55_w143, c0_n55_w144, c0_n55_w145, c0_n55_w146, c0_n55_w147, c0_n55_w148, c0_n55_w149, c0_n55_w150, c0_n55_w151, c0_n55_w152, c0_n55_w153, c0_n55_w154, c0_n55_w155, c0_n55_w156, c0_n55_w157, c0_n55_w158, c0_n55_w159, c0_n55_w160, c0_n55_w161, c0_n55_w162, c0_n55_w163, c0_n55_w164, c0_n55_w165, c0_n55_w166, c0_n55_w167, c0_n55_w168, c0_n55_w169, c0_n55_w170, c0_n55_w171, c0_n55_w172, c0_n55_w173, c0_n55_w174, c0_n55_w175, c0_n55_w176, c0_n55_w177, c0_n55_w178, c0_n55_w179, c0_n55_w180, c0_n55_w181, c0_n55_w182, c0_n55_w183, c0_n55_w184, c0_n55_w185, c0_n55_w186, c0_n55_w187, c0_n55_w188, c0_n55_w189, c0_n55_w190, c0_n55_w191, c0_n55_w192, c0_n55_w193, c0_n55_w194, c0_n55_w195, c0_n55_w196, c0_n55_w197, c0_n55_w198, c0_n55_w199, c0_n55_w200, c0_n56_w1, c0_n56_w2, c0_n56_w3, c0_n56_w4, c0_n56_w5, c0_n56_w6, c0_n56_w7, c0_n56_w8, c0_n56_w9, c0_n56_w10, c0_n56_w11, c0_n56_w12, c0_n56_w13, c0_n56_w14, c0_n56_w15, c0_n56_w16, c0_n56_w17, c0_n56_w18, c0_n56_w19, c0_n56_w20, c0_n56_w21, c0_n56_w22, c0_n56_w23, c0_n56_w24, c0_n56_w25, c0_n56_w26, c0_n56_w27, c0_n56_w28, c0_n56_w29, c0_n56_w30, c0_n56_w31, c0_n56_w32, c0_n56_w33, c0_n56_w34, c0_n56_w35, c0_n56_w36, c0_n56_w37, c0_n56_w38, c0_n56_w39, c0_n56_w40, c0_n56_w41, c0_n56_w42, c0_n56_w43, c0_n56_w44, c0_n56_w45, c0_n56_w46, c0_n56_w47, c0_n56_w48, c0_n56_w49, c0_n56_w50, c0_n56_w51, c0_n56_w52, c0_n56_w53, c0_n56_w54, c0_n56_w55, c0_n56_w56, c0_n56_w57, c0_n56_w58, c0_n56_w59, c0_n56_w60, c0_n56_w61, c0_n56_w62, c0_n56_w63, c0_n56_w64, c0_n56_w65, c0_n56_w66, c0_n56_w67, c0_n56_w68, c0_n56_w69, c0_n56_w70, c0_n56_w71, c0_n56_w72, c0_n56_w73, c0_n56_w74, c0_n56_w75, c0_n56_w76, c0_n56_w77, c0_n56_w78, c0_n56_w79, c0_n56_w80, c0_n56_w81, c0_n56_w82, c0_n56_w83, c0_n56_w84, c0_n56_w85, c0_n56_w86, c0_n56_w87, c0_n56_w88, c0_n56_w89, c0_n56_w90, c0_n56_w91, c0_n56_w92, c0_n56_w93, c0_n56_w94, c0_n56_w95, c0_n56_w96, c0_n56_w97, c0_n56_w98, c0_n56_w99, c0_n56_w100, c0_n56_w101, c0_n56_w102, c0_n56_w103, c0_n56_w104, c0_n56_w105, c0_n56_w106, c0_n56_w107, c0_n56_w108, c0_n56_w109, c0_n56_w110, c0_n56_w111, c0_n56_w112, c0_n56_w113, c0_n56_w114, c0_n56_w115, c0_n56_w116, c0_n56_w117, c0_n56_w118, c0_n56_w119, c0_n56_w120, c0_n56_w121, c0_n56_w122, c0_n56_w123, c0_n56_w124, c0_n56_w125, c0_n56_w126, c0_n56_w127, c0_n56_w128, c0_n56_w129, c0_n56_w130, c0_n56_w131, c0_n56_w132, c0_n56_w133, c0_n56_w134, c0_n56_w135, c0_n56_w136, c0_n56_w137, c0_n56_w138, c0_n56_w139, c0_n56_w140, c0_n56_w141, c0_n56_w142, c0_n56_w143, c0_n56_w144, c0_n56_w145, c0_n56_w146, c0_n56_w147, c0_n56_w148, c0_n56_w149, c0_n56_w150, c0_n56_w151, c0_n56_w152, c0_n56_w153, c0_n56_w154, c0_n56_w155, c0_n56_w156, c0_n56_w157, c0_n56_w158, c0_n56_w159, c0_n56_w160, c0_n56_w161, c0_n56_w162, c0_n56_w163, c0_n56_w164, c0_n56_w165, c0_n56_w166, c0_n56_w167, c0_n56_w168, c0_n56_w169, c0_n56_w170, c0_n56_w171, c0_n56_w172, c0_n56_w173, c0_n56_w174, c0_n56_w175, c0_n56_w176, c0_n56_w177, c0_n56_w178, c0_n56_w179, c0_n56_w180, c0_n56_w181, c0_n56_w182, c0_n56_w183, c0_n56_w184, c0_n56_w185, c0_n56_w186, c0_n56_w187, c0_n56_w188, c0_n56_w189, c0_n56_w190, c0_n56_w191, c0_n56_w192, c0_n56_w193, c0_n56_w194, c0_n56_w195, c0_n56_w196, c0_n56_w197, c0_n56_w198, c0_n56_w199, c0_n56_w200, c0_n57_w1, c0_n57_w2, c0_n57_w3, c0_n57_w4, c0_n57_w5, c0_n57_w6, c0_n57_w7, c0_n57_w8, c0_n57_w9, c0_n57_w10, c0_n57_w11, c0_n57_w12, c0_n57_w13, c0_n57_w14, c0_n57_w15, c0_n57_w16, c0_n57_w17, c0_n57_w18, c0_n57_w19, c0_n57_w20, c0_n57_w21, c0_n57_w22, c0_n57_w23, c0_n57_w24, c0_n57_w25, c0_n57_w26, c0_n57_w27, c0_n57_w28, c0_n57_w29, c0_n57_w30, c0_n57_w31, c0_n57_w32, c0_n57_w33, c0_n57_w34, c0_n57_w35, c0_n57_w36, c0_n57_w37, c0_n57_w38, c0_n57_w39, c0_n57_w40, c0_n57_w41, c0_n57_w42, c0_n57_w43, c0_n57_w44, c0_n57_w45, c0_n57_w46, c0_n57_w47, c0_n57_w48, c0_n57_w49, c0_n57_w50, c0_n57_w51, c0_n57_w52, c0_n57_w53, c0_n57_w54, c0_n57_w55, c0_n57_w56, c0_n57_w57, c0_n57_w58, c0_n57_w59, c0_n57_w60, c0_n57_w61, c0_n57_w62, c0_n57_w63, c0_n57_w64, c0_n57_w65, c0_n57_w66, c0_n57_w67, c0_n57_w68, c0_n57_w69, c0_n57_w70, c0_n57_w71, c0_n57_w72, c0_n57_w73, c0_n57_w74, c0_n57_w75, c0_n57_w76, c0_n57_w77, c0_n57_w78, c0_n57_w79, c0_n57_w80, c0_n57_w81, c0_n57_w82, c0_n57_w83, c0_n57_w84, c0_n57_w85, c0_n57_w86, c0_n57_w87, c0_n57_w88, c0_n57_w89, c0_n57_w90, c0_n57_w91, c0_n57_w92, c0_n57_w93, c0_n57_w94, c0_n57_w95, c0_n57_w96, c0_n57_w97, c0_n57_w98, c0_n57_w99, c0_n57_w100, c0_n57_w101, c0_n57_w102, c0_n57_w103, c0_n57_w104, c0_n57_w105, c0_n57_w106, c0_n57_w107, c0_n57_w108, c0_n57_w109, c0_n57_w110, c0_n57_w111, c0_n57_w112, c0_n57_w113, c0_n57_w114, c0_n57_w115, c0_n57_w116, c0_n57_w117, c0_n57_w118, c0_n57_w119, c0_n57_w120, c0_n57_w121, c0_n57_w122, c0_n57_w123, c0_n57_w124, c0_n57_w125, c0_n57_w126, c0_n57_w127, c0_n57_w128, c0_n57_w129, c0_n57_w130, c0_n57_w131, c0_n57_w132, c0_n57_w133, c0_n57_w134, c0_n57_w135, c0_n57_w136, c0_n57_w137, c0_n57_w138, c0_n57_w139, c0_n57_w140, c0_n57_w141, c0_n57_w142, c0_n57_w143, c0_n57_w144, c0_n57_w145, c0_n57_w146, c0_n57_w147, c0_n57_w148, c0_n57_w149, c0_n57_w150, c0_n57_w151, c0_n57_w152, c0_n57_w153, c0_n57_w154, c0_n57_w155, c0_n57_w156, c0_n57_w157, c0_n57_w158, c0_n57_w159, c0_n57_w160, c0_n57_w161, c0_n57_w162, c0_n57_w163, c0_n57_w164, c0_n57_w165, c0_n57_w166, c0_n57_w167, c0_n57_w168, c0_n57_w169, c0_n57_w170, c0_n57_w171, c0_n57_w172, c0_n57_w173, c0_n57_w174, c0_n57_w175, c0_n57_w176, c0_n57_w177, c0_n57_w178, c0_n57_w179, c0_n57_w180, c0_n57_w181, c0_n57_w182, c0_n57_w183, c0_n57_w184, c0_n57_w185, c0_n57_w186, c0_n57_w187, c0_n57_w188, c0_n57_w189, c0_n57_w190, c0_n57_w191, c0_n57_w192, c0_n57_w193, c0_n57_w194, c0_n57_w195, c0_n57_w196, c0_n57_w197, c0_n57_w198, c0_n57_w199, c0_n57_w200, c0_n58_w1, c0_n58_w2, c0_n58_w3, c0_n58_w4, c0_n58_w5, c0_n58_w6, c0_n58_w7, c0_n58_w8, c0_n58_w9, c0_n58_w10, c0_n58_w11, c0_n58_w12, c0_n58_w13, c0_n58_w14, c0_n58_w15, c0_n58_w16, c0_n58_w17, c0_n58_w18, c0_n58_w19, c0_n58_w20, c0_n58_w21, c0_n58_w22, c0_n58_w23, c0_n58_w24, c0_n58_w25, c0_n58_w26, c0_n58_w27, c0_n58_w28, c0_n58_w29, c0_n58_w30, c0_n58_w31, c0_n58_w32, c0_n58_w33, c0_n58_w34, c0_n58_w35, c0_n58_w36, c0_n58_w37, c0_n58_w38, c0_n58_w39, c0_n58_w40, c0_n58_w41, c0_n58_w42, c0_n58_w43, c0_n58_w44, c0_n58_w45, c0_n58_w46, c0_n58_w47, c0_n58_w48, c0_n58_w49, c0_n58_w50, c0_n58_w51, c0_n58_w52, c0_n58_w53, c0_n58_w54, c0_n58_w55, c0_n58_w56, c0_n58_w57, c0_n58_w58, c0_n58_w59, c0_n58_w60, c0_n58_w61, c0_n58_w62, c0_n58_w63, c0_n58_w64, c0_n58_w65, c0_n58_w66, c0_n58_w67, c0_n58_w68, c0_n58_w69, c0_n58_w70, c0_n58_w71, c0_n58_w72, c0_n58_w73, c0_n58_w74, c0_n58_w75, c0_n58_w76, c0_n58_w77, c0_n58_w78, c0_n58_w79, c0_n58_w80, c0_n58_w81, c0_n58_w82, c0_n58_w83, c0_n58_w84, c0_n58_w85, c0_n58_w86, c0_n58_w87, c0_n58_w88, c0_n58_w89, c0_n58_w90, c0_n58_w91, c0_n58_w92, c0_n58_w93, c0_n58_w94, c0_n58_w95, c0_n58_w96, c0_n58_w97, c0_n58_w98, c0_n58_w99, c0_n58_w100, c0_n58_w101, c0_n58_w102, c0_n58_w103, c0_n58_w104, c0_n58_w105, c0_n58_w106, c0_n58_w107, c0_n58_w108, c0_n58_w109, c0_n58_w110, c0_n58_w111, c0_n58_w112, c0_n58_w113, c0_n58_w114, c0_n58_w115, c0_n58_w116, c0_n58_w117, c0_n58_w118, c0_n58_w119, c0_n58_w120, c0_n58_w121, c0_n58_w122, c0_n58_w123, c0_n58_w124, c0_n58_w125, c0_n58_w126, c0_n58_w127, c0_n58_w128, c0_n58_w129, c0_n58_w130, c0_n58_w131, c0_n58_w132, c0_n58_w133, c0_n58_w134, c0_n58_w135, c0_n58_w136, c0_n58_w137, c0_n58_w138, c0_n58_w139, c0_n58_w140, c0_n58_w141, c0_n58_w142, c0_n58_w143, c0_n58_w144, c0_n58_w145, c0_n58_w146, c0_n58_w147, c0_n58_w148, c0_n58_w149, c0_n58_w150, c0_n58_w151, c0_n58_w152, c0_n58_w153, c0_n58_w154, c0_n58_w155, c0_n58_w156, c0_n58_w157, c0_n58_w158, c0_n58_w159, c0_n58_w160, c0_n58_w161, c0_n58_w162, c0_n58_w163, c0_n58_w164, c0_n58_w165, c0_n58_w166, c0_n58_w167, c0_n58_w168, c0_n58_w169, c0_n58_w170, c0_n58_w171, c0_n58_w172, c0_n58_w173, c0_n58_w174, c0_n58_w175, c0_n58_w176, c0_n58_w177, c0_n58_w178, c0_n58_w179, c0_n58_w180, c0_n58_w181, c0_n58_w182, c0_n58_w183, c0_n58_w184, c0_n58_w185, c0_n58_w186, c0_n58_w187, c0_n58_w188, c0_n58_w189, c0_n58_w190, c0_n58_w191, c0_n58_w192, c0_n58_w193, c0_n58_w194, c0_n58_w195, c0_n58_w196, c0_n58_w197, c0_n58_w198, c0_n58_w199, c0_n58_w200, c0_n59_w1, c0_n59_w2, c0_n59_w3, c0_n59_w4, c0_n59_w5, c0_n59_w6, c0_n59_w7, c0_n59_w8, c0_n59_w9, c0_n59_w10, c0_n59_w11, c0_n59_w12, c0_n59_w13, c0_n59_w14, c0_n59_w15, c0_n59_w16, c0_n59_w17, c0_n59_w18, c0_n59_w19, c0_n59_w20, c0_n59_w21, c0_n59_w22, c0_n59_w23, c0_n59_w24, c0_n59_w25, c0_n59_w26, c0_n59_w27, c0_n59_w28, c0_n59_w29, c0_n59_w30, c0_n59_w31, c0_n59_w32, c0_n59_w33, c0_n59_w34, c0_n59_w35, c0_n59_w36, c0_n59_w37, c0_n59_w38, c0_n59_w39, c0_n59_w40, c0_n59_w41, c0_n59_w42, c0_n59_w43, c0_n59_w44, c0_n59_w45, c0_n59_w46, c0_n59_w47, c0_n59_w48, c0_n59_w49, c0_n59_w50, c0_n59_w51, c0_n59_w52, c0_n59_w53, c0_n59_w54, c0_n59_w55, c0_n59_w56, c0_n59_w57, c0_n59_w58, c0_n59_w59, c0_n59_w60, c0_n59_w61, c0_n59_w62, c0_n59_w63, c0_n59_w64, c0_n59_w65, c0_n59_w66, c0_n59_w67, c0_n59_w68, c0_n59_w69, c0_n59_w70, c0_n59_w71, c0_n59_w72, c0_n59_w73, c0_n59_w74, c0_n59_w75, c0_n59_w76, c0_n59_w77, c0_n59_w78, c0_n59_w79, c0_n59_w80, c0_n59_w81, c0_n59_w82, c0_n59_w83, c0_n59_w84, c0_n59_w85, c0_n59_w86, c0_n59_w87, c0_n59_w88, c0_n59_w89, c0_n59_w90, c0_n59_w91, c0_n59_w92, c0_n59_w93, c0_n59_w94, c0_n59_w95, c0_n59_w96, c0_n59_w97, c0_n59_w98, c0_n59_w99, c0_n59_w100, c0_n59_w101, c0_n59_w102, c0_n59_w103, c0_n59_w104, c0_n59_w105, c0_n59_w106, c0_n59_w107, c0_n59_w108, c0_n59_w109, c0_n59_w110, c0_n59_w111, c0_n59_w112, c0_n59_w113, c0_n59_w114, c0_n59_w115, c0_n59_w116, c0_n59_w117, c0_n59_w118, c0_n59_w119, c0_n59_w120, c0_n59_w121, c0_n59_w122, c0_n59_w123, c0_n59_w124, c0_n59_w125, c0_n59_w126, c0_n59_w127, c0_n59_w128, c0_n59_w129, c0_n59_w130, c0_n59_w131, c0_n59_w132, c0_n59_w133, c0_n59_w134, c0_n59_w135, c0_n59_w136, c0_n59_w137, c0_n59_w138, c0_n59_w139, c0_n59_w140, c0_n59_w141, c0_n59_w142, c0_n59_w143, c0_n59_w144, c0_n59_w145, c0_n59_w146, c0_n59_w147, c0_n59_w148, c0_n59_w149, c0_n59_w150, c0_n59_w151, c0_n59_w152, c0_n59_w153, c0_n59_w154, c0_n59_w155, c0_n59_w156, c0_n59_w157, c0_n59_w158, c0_n59_w159, c0_n59_w160, c0_n59_w161, c0_n59_w162, c0_n59_w163, c0_n59_w164, c0_n59_w165, c0_n59_w166, c0_n59_w167, c0_n59_w168, c0_n59_w169, c0_n59_w170, c0_n59_w171, c0_n59_w172, c0_n59_w173, c0_n59_w174, c0_n59_w175, c0_n59_w176, c0_n59_w177, c0_n59_w178, c0_n59_w179, c0_n59_w180, c0_n59_w181, c0_n59_w182, c0_n59_w183, c0_n59_w184, c0_n59_w185, c0_n59_w186, c0_n59_w187, c0_n59_w188, c0_n59_w189, c0_n59_w190, c0_n59_w191, c0_n59_w192, c0_n59_w193, c0_n59_w194, c0_n59_w195, c0_n59_w196, c0_n59_w197, c0_n59_w198, c0_n59_w199, c0_n59_w200, c0_n60_w1, c0_n60_w2, c0_n60_w3, c0_n60_w4, c0_n60_w5, c0_n60_w6, c0_n60_w7, c0_n60_w8, c0_n60_w9, c0_n60_w10, c0_n60_w11, c0_n60_w12, c0_n60_w13, c0_n60_w14, c0_n60_w15, c0_n60_w16, c0_n60_w17, c0_n60_w18, c0_n60_w19, c0_n60_w20, c0_n60_w21, c0_n60_w22, c0_n60_w23, c0_n60_w24, c0_n60_w25, c0_n60_w26, c0_n60_w27, c0_n60_w28, c0_n60_w29, c0_n60_w30, c0_n60_w31, c0_n60_w32, c0_n60_w33, c0_n60_w34, c0_n60_w35, c0_n60_w36, c0_n60_w37, c0_n60_w38, c0_n60_w39, c0_n60_w40, c0_n60_w41, c0_n60_w42, c0_n60_w43, c0_n60_w44, c0_n60_w45, c0_n60_w46, c0_n60_w47, c0_n60_w48, c0_n60_w49, c0_n60_w50, c0_n60_w51, c0_n60_w52, c0_n60_w53, c0_n60_w54, c0_n60_w55, c0_n60_w56, c0_n60_w57, c0_n60_w58, c0_n60_w59, c0_n60_w60, c0_n60_w61, c0_n60_w62, c0_n60_w63, c0_n60_w64, c0_n60_w65, c0_n60_w66, c0_n60_w67, c0_n60_w68, c0_n60_w69, c0_n60_w70, c0_n60_w71, c0_n60_w72, c0_n60_w73, c0_n60_w74, c0_n60_w75, c0_n60_w76, c0_n60_w77, c0_n60_w78, c0_n60_w79, c0_n60_w80, c0_n60_w81, c0_n60_w82, c0_n60_w83, c0_n60_w84, c0_n60_w85, c0_n60_w86, c0_n60_w87, c0_n60_w88, c0_n60_w89, c0_n60_w90, c0_n60_w91, c0_n60_w92, c0_n60_w93, c0_n60_w94, c0_n60_w95, c0_n60_w96, c0_n60_w97, c0_n60_w98, c0_n60_w99, c0_n60_w100, c0_n60_w101, c0_n60_w102, c0_n60_w103, c0_n60_w104, c0_n60_w105, c0_n60_w106, c0_n60_w107, c0_n60_w108, c0_n60_w109, c0_n60_w110, c0_n60_w111, c0_n60_w112, c0_n60_w113, c0_n60_w114, c0_n60_w115, c0_n60_w116, c0_n60_w117, c0_n60_w118, c0_n60_w119, c0_n60_w120, c0_n60_w121, c0_n60_w122, c0_n60_w123, c0_n60_w124, c0_n60_w125, c0_n60_w126, c0_n60_w127, c0_n60_w128, c0_n60_w129, c0_n60_w130, c0_n60_w131, c0_n60_w132, c0_n60_w133, c0_n60_w134, c0_n60_w135, c0_n60_w136, c0_n60_w137, c0_n60_w138, c0_n60_w139, c0_n60_w140, c0_n60_w141, c0_n60_w142, c0_n60_w143, c0_n60_w144, c0_n60_w145, c0_n60_w146, c0_n60_w147, c0_n60_w148, c0_n60_w149, c0_n60_w150, c0_n60_w151, c0_n60_w152, c0_n60_w153, c0_n60_w154, c0_n60_w155, c0_n60_w156, c0_n60_w157, c0_n60_w158, c0_n60_w159, c0_n60_w160, c0_n60_w161, c0_n60_w162, c0_n60_w163, c0_n60_w164, c0_n60_w165, c0_n60_w166, c0_n60_w167, c0_n60_w168, c0_n60_w169, c0_n60_w170, c0_n60_w171, c0_n60_w172, c0_n60_w173, c0_n60_w174, c0_n60_w175, c0_n60_w176, c0_n60_w177, c0_n60_w178, c0_n60_w179, c0_n60_w180, c0_n60_w181, c0_n60_w182, c0_n60_w183, c0_n60_w184, c0_n60_w185, c0_n60_w186, c0_n60_w187, c0_n60_w188, c0_n60_w189, c0_n60_w190, c0_n60_w191, c0_n60_w192, c0_n60_w193, c0_n60_w194, c0_n60_w195, c0_n60_w196, c0_n60_w197, c0_n60_w198, c0_n60_w199, c0_n60_w200, c0_n61_w1, c0_n61_w2, c0_n61_w3, c0_n61_w4, c0_n61_w5, c0_n61_w6, c0_n61_w7, c0_n61_w8, c0_n61_w9, c0_n61_w10, c0_n61_w11, c0_n61_w12, c0_n61_w13, c0_n61_w14, c0_n61_w15, c0_n61_w16, c0_n61_w17, c0_n61_w18, c0_n61_w19, c0_n61_w20, c0_n61_w21, c0_n61_w22, c0_n61_w23, c0_n61_w24, c0_n61_w25, c0_n61_w26, c0_n61_w27, c0_n61_w28, c0_n61_w29, c0_n61_w30, c0_n61_w31, c0_n61_w32, c0_n61_w33, c0_n61_w34, c0_n61_w35, c0_n61_w36, c0_n61_w37, c0_n61_w38, c0_n61_w39, c0_n61_w40, c0_n61_w41, c0_n61_w42, c0_n61_w43, c0_n61_w44, c0_n61_w45, c0_n61_w46, c0_n61_w47, c0_n61_w48, c0_n61_w49, c0_n61_w50, c0_n61_w51, c0_n61_w52, c0_n61_w53, c0_n61_w54, c0_n61_w55, c0_n61_w56, c0_n61_w57, c0_n61_w58, c0_n61_w59, c0_n61_w60, c0_n61_w61, c0_n61_w62, c0_n61_w63, c0_n61_w64, c0_n61_w65, c0_n61_w66, c0_n61_w67, c0_n61_w68, c0_n61_w69, c0_n61_w70, c0_n61_w71, c0_n61_w72, c0_n61_w73, c0_n61_w74, c0_n61_w75, c0_n61_w76, c0_n61_w77, c0_n61_w78, c0_n61_w79, c0_n61_w80, c0_n61_w81, c0_n61_w82, c0_n61_w83, c0_n61_w84, c0_n61_w85, c0_n61_w86, c0_n61_w87, c0_n61_w88, c0_n61_w89, c0_n61_w90, c0_n61_w91, c0_n61_w92, c0_n61_w93, c0_n61_w94, c0_n61_w95, c0_n61_w96, c0_n61_w97, c0_n61_w98, c0_n61_w99, c0_n61_w100, c0_n61_w101, c0_n61_w102, c0_n61_w103, c0_n61_w104, c0_n61_w105, c0_n61_w106, c0_n61_w107, c0_n61_w108, c0_n61_w109, c0_n61_w110, c0_n61_w111, c0_n61_w112, c0_n61_w113, c0_n61_w114, c0_n61_w115, c0_n61_w116, c0_n61_w117, c0_n61_w118, c0_n61_w119, c0_n61_w120, c0_n61_w121, c0_n61_w122, c0_n61_w123, c0_n61_w124, c0_n61_w125, c0_n61_w126, c0_n61_w127, c0_n61_w128, c0_n61_w129, c0_n61_w130, c0_n61_w131, c0_n61_w132, c0_n61_w133, c0_n61_w134, c0_n61_w135, c0_n61_w136, c0_n61_w137, c0_n61_w138, c0_n61_w139, c0_n61_w140, c0_n61_w141, c0_n61_w142, c0_n61_w143, c0_n61_w144, c0_n61_w145, c0_n61_w146, c0_n61_w147, c0_n61_w148, c0_n61_w149, c0_n61_w150, c0_n61_w151, c0_n61_w152, c0_n61_w153, c0_n61_w154, c0_n61_w155, c0_n61_w156, c0_n61_w157, c0_n61_w158, c0_n61_w159, c0_n61_w160, c0_n61_w161, c0_n61_w162, c0_n61_w163, c0_n61_w164, c0_n61_w165, c0_n61_w166, c0_n61_w167, c0_n61_w168, c0_n61_w169, c0_n61_w170, c0_n61_w171, c0_n61_w172, c0_n61_w173, c0_n61_w174, c0_n61_w175, c0_n61_w176, c0_n61_w177, c0_n61_w178, c0_n61_w179, c0_n61_w180, c0_n61_w181, c0_n61_w182, c0_n61_w183, c0_n61_w184, c0_n61_w185, c0_n61_w186, c0_n61_w187, c0_n61_w188, c0_n61_w189, c0_n61_w190, c0_n61_w191, c0_n61_w192, c0_n61_w193, c0_n61_w194, c0_n61_w195, c0_n61_w196, c0_n61_w197, c0_n61_w198, c0_n61_w199, c0_n61_w200, c0_n62_w1, c0_n62_w2, c0_n62_w3, c0_n62_w4, c0_n62_w5, c0_n62_w6, c0_n62_w7, c0_n62_w8, c0_n62_w9, c0_n62_w10, c0_n62_w11, c0_n62_w12, c0_n62_w13, c0_n62_w14, c0_n62_w15, c0_n62_w16, c0_n62_w17, c0_n62_w18, c0_n62_w19, c0_n62_w20, c0_n62_w21, c0_n62_w22, c0_n62_w23, c0_n62_w24, c0_n62_w25, c0_n62_w26, c0_n62_w27, c0_n62_w28, c0_n62_w29, c0_n62_w30, c0_n62_w31, c0_n62_w32, c0_n62_w33, c0_n62_w34, c0_n62_w35, c0_n62_w36, c0_n62_w37, c0_n62_w38, c0_n62_w39, c0_n62_w40, c0_n62_w41, c0_n62_w42, c0_n62_w43, c0_n62_w44, c0_n62_w45, c0_n62_w46, c0_n62_w47, c0_n62_w48, c0_n62_w49, c0_n62_w50, c0_n62_w51, c0_n62_w52, c0_n62_w53, c0_n62_w54, c0_n62_w55, c0_n62_w56, c0_n62_w57, c0_n62_w58, c0_n62_w59, c0_n62_w60, c0_n62_w61, c0_n62_w62, c0_n62_w63, c0_n62_w64, c0_n62_w65, c0_n62_w66, c0_n62_w67, c0_n62_w68, c0_n62_w69, c0_n62_w70, c0_n62_w71, c0_n62_w72, c0_n62_w73, c0_n62_w74, c0_n62_w75, c0_n62_w76, c0_n62_w77, c0_n62_w78, c0_n62_w79, c0_n62_w80, c0_n62_w81, c0_n62_w82, c0_n62_w83, c0_n62_w84, c0_n62_w85, c0_n62_w86, c0_n62_w87, c0_n62_w88, c0_n62_w89, c0_n62_w90, c0_n62_w91, c0_n62_w92, c0_n62_w93, c0_n62_w94, c0_n62_w95, c0_n62_w96, c0_n62_w97, c0_n62_w98, c0_n62_w99, c0_n62_w100, c0_n62_w101, c0_n62_w102, c0_n62_w103, c0_n62_w104, c0_n62_w105, c0_n62_w106, c0_n62_w107, c0_n62_w108, c0_n62_w109, c0_n62_w110, c0_n62_w111, c0_n62_w112, c0_n62_w113, c0_n62_w114, c0_n62_w115, c0_n62_w116, c0_n62_w117, c0_n62_w118, c0_n62_w119, c0_n62_w120, c0_n62_w121, c0_n62_w122, c0_n62_w123, c0_n62_w124, c0_n62_w125, c0_n62_w126, c0_n62_w127, c0_n62_w128, c0_n62_w129, c0_n62_w130, c0_n62_w131, c0_n62_w132, c0_n62_w133, c0_n62_w134, c0_n62_w135, c0_n62_w136, c0_n62_w137, c0_n62_w138, c0_n62_w139, c0_n62_w140, c0_n62_w141, c0_n62_w142, c0_n62_w143, c0_n62_w144, c0_n62_w145, c0_n62_w146, c0_n62_w147, c0_n62_w148, c0_n62_w149, c0_n62_w150, c0_n62_w151, c0_n62_w152, c0_n62_w153, c0_n62_w154, c0_n62_w155, c0_n62_w156, c0_n62_w157, c0_n62_w158, c0_n62_w159, c0_n62_w160, c0_n62_w161, c0_n62_w162, c0_n62_w163, c0_n62_w164, c0_n62_w165, c0_n62_w166, c0_n62_w167, c0_n62_w168, c0_n62_w169, c0_n62_w170, c0_n62_w171, c0_n62_w172, c0_n62_w173, c0_n62_w174, c0_n62_w175, c0_n62_w176, c0_n62_w177, c0_n62_w178, c0_n62_w179, c0_n62_w180, c0_n62_w181, c0_n62_w182, c0_n62_w183, c0_n62_w184, c0_n62_w185, c0_n62_w186, c0_n62_w187, c0_n62_w188, c0_n62_w189, c0_n62_w190, c0_n62_w191, c0_n62_w192, c0_n62_w193, c0_n62_w194, c0_n62_w195, c0_n62_w196, c0_n62_w197, c0_n62_w198, c0_n62_w199, c0_n62_w200, c0_n63_w1, c0_n63_w2, c0_n63_w3, c0_n63_w4, c0_n63_w5, c0_n63_w6, c0_n63_w7, c0_n63_w8, c0_n63_w9, c0_n63_w10, c0_n63_w11, c0_n63_w12, c0_n63_w13, c0_n63_w14, c0_n63_w15, c0_n63_w16, c0_n63_w17, c0_n63_w18, c0_n63_w19, c0_n63_w20, c0_n63_w21, c0_n63_w22, c0_n63_w23, c0_n63_w24, c0_n63_w25, c0_n63_w26, c0_n63_w27, c0_n63_w28, c0_n63_w29, c0_n63_w30, c0_n63_w31, c0_n63_w32, c0_n63_w33, c0_n63_w34, c0_n63_w35, c0_n63_w36, c0_n63_w37, c0_n63_w38, c0_n63_w39, c0_n63_w40, c0_n63_w41, c0_n63_w42, c0_n63_w43, c0_n63_w44, c0_n63_w45, c0_n63_w46, c0_n63_w47, c0_n63_w48, c0_n63_w49, c0_n63_w50, c0_n63_w51, c0_n63_w52, c0_n63_w53, c0_n63_w54, c0_n63_w55, c0_n63_w56, c0_n63_w57, c0_n63_w58, c0_n63_w59, c0_n63_w60, c0_n63_w61, c0_n63_w62, c0_n63_w63, c0_n63_w64, c0_n63_w65, c0_n63_w66, c0_n63_w67, c0_n63_w68, c0_n63_w69, c0_n63_w70, c0_n63_w71, c0_n63_w72, c0_n63_w73, c0_n63_w74, c0_n63_w75, c0_n63_w76, c0_n63_w77, c0_n63_w78, c0_n63_w79, c0_n63_w80, c0_n63_w81, c0_n63_w82, c0_n63_w83, c0_n63_w84, c0_n63_w85, c0_n63_w86, c0_n63_w87, c0_n63_w88, c0_n63_w89, c0_n63_w90, c0_n63_w91, c0_n63_w92, c0_n63_w93, c0_n63_w94, c0_n63_w95, c0_n63_w96, c0_n63_w97, c0_n63_w98, c0_n63_w99, c0_n63_w100, c0_n63_w101, c0_n63_w102, c0_n63_w103, c0_n63_w104, c0_n63_w105, c0_n63_w106, c0_n63_w107, c0_n63_w108, c0_n63_w109, c0_n63_w110, c0_n63_w111, c0_n63_w112, c0_n63_w113, c0_n63_w114, c0_n63_w115, c0_n63_w116, c0_n63_w117, c0_n63_w118, c0_n63_w119, c0_n63_w120, c0_n63_w121, c0_n63_w122, c0_n63_w123, c0_n63_w124, c0_n63_w125, c0_n63_w126, c0_n63_w127, c0_n63_w128, c0_n63_w129, c0_n63_w130, c0_n63_w131, c0_n63_w132, c0_n63_w133, c0_n63_w134, c0_n63_w135, c0_n63_w136, c0_n63_w137, c0_n63_w138, c0_n63_w139, c0_n63_w140, c0_n63_w141, c0_n63_w142, c0_n63_w143, c0_n63_w144, c0_n63_w145, c0_n63_w146, c0_n63_w147, c0_n63_w148, c0_n63_w149, c0_n63_w150, c0_n63_w151, c0_n63_w152, c0_n63_w153, c0_n63_w154, c0_n63_w155, c0_n63_w156, c0_n63_w157, c0_n63_w158, c0_n63_w159, c0_n63_w160, c0_n63_w161, c0_n63_w162, c0_n63_w163, c0_n63_w164, c0_n63_w165, c0_n63_w166, c0_n63_w167, c0_n63_w168, c0_n63_w169, c0_n63_w170, c0_n63_w171, c0_n63_w172, c0_n63_w173, c0_n63_w174, c0_n63_w175, c0_n63_w176, c0_n63_w177, c0_n63_w178, c0_n63_w179, c0_n63_w180, c0_n63_w181, c0_n63_w182, c0_n63_w183, c0_n63_w184, c0_n63_w185, c0_n63_w186, c0_n63_w187, c0_n63_w188, c0_n63_w189, c0_n63_w190, c0_n63_w191, c0_n63_w192, c0_n63_w193, c0_n63_w194, c0_n63_w195, c0_n63_w196, c0_n63_w197, c0_n63_w198, c0_n63_w199, c0_n63_w200, c0_n64_w1, c0_n64_w2, c0_n64_w3, c0_n64_w4, c0_n64_w5, c0_n64_w6, c0_n64_w7, c0_n64_w8, c0_n64_w9, c0_n64_w10, c0_n64_w11, c0_n64_w12, c0_n64_w13, c0_n64_w14, c0_n64_w15, c0_n64_w16, c0_n64_w17, c0_n64_w18, c0_n64_w19, c0_n64_w20, c0_n64_w21, c0_n64_w22, c0_n64_w23, c0_n64_w24, c0_n64_w25, c0_n64_w26, c0_n64_w27, c0_n64_w28, c0_n64_w29, c0_n64_w30, c0_n64_w31, c0_n64_w32, c0_n64_w33, c0_n64_w34, c0_n64_w35, c0_n64_w36, c0_n64_w37, c0_n64_w38, c0_n64_w39, c0_n64_w40, c0_n64_w41, c0_n64_w42, c0_n64_w43, c0_n64_w44, c0_n64_w45, c0_n64_w46, c0_n64_w47, c0_n64_w48, c0_n64_w49, c0_n64_w50, c0_n64_w51, c0_n64_w52, c0_n64_w53, c0_n64_w54, c0_n64_w55, c0_n64_w56, c0_n64_w57, c0_n64_w58, c0_n64_w59, c0_n64_w60, c0_n64_w61, c0_n64_w62, c0_n64_w63, c0_n64_w64, c0_n64_w65, c0_n64_w66, c0_n64_w67, c0_n64_w68, c0_n64_w69, c0_n64_w70, c0_n64_w71, c0_n64_w72, c0_n64_w73, c0_n64_w74, c0_n64_w75, c0_n64_w76, c0_n64_w77, c0_n64_w78, c0_n64_w79, c0_n64_w80, c0_n64_w81, c0_n64_w82, c0_n64_w83, c0_n64_w84, c0_n64_w85, c0_n64_w86, c0_n64_w87, c0_n64_w88, c0_n64_w89, c0_n64_w90, c0_n64_w91, c0_n64_w92, c0_n64_w93, c0_n64_w94, c0_n64_w95, c0_n64_w96, c0_n64_w97, c0_n64_w98, c0_n64_w99, c0_n64_w100, c0_n64_w101, c0_n64_w102, c0_n64_w103, c0_n64_w104, c0_n64_w105, c0_n64_w106, c0_n64_w107, c0_n64_w108, c0_n64_w109, c0_n64_w110, c0_n64_w111, c0_n64_w112, c0_n64_w113, c0_n64_w114, c0_n64_w115, c0_n64_w116, c0_n64_w117, c0_n64_w118, c0_n64_w119, c0_n64_w120, c0_n64_w121, c0_n64_w122, c0_n64_w123, c0_n64_w124, c0_n64_w125, c0_n64_w126, c0_n64_w127, c0_n64_w128, c0_n64_w129, c0_n64_w130, c0_n64_w131, c0_n64_w132, c0_n64_w133, c0_n64_w134, c0_n64_w135, c0_n64_w136, c0_n64_w137, c0_n64_w138, c0_n64_w139, c0_n64_w140, c0_n64_w141, c0_n64_w142, c0_n64_w143, c0_n64_w144, c0_n64_w145, c0_n64_w146, c0_n64_w147, c0_n64_w148, c0_n64_w149, c0_n64_w150, c0_n64_w151, c0_n64_w152, c0_n64_w153, c0_n64_w154, c0_n64_w155, c0_n64_w156, c0_n64_w157, c0_n64_w158, c0_n64_w159, c0_n64_w160, c0_n64_w161, c0_n64_w162, c0_n64_w163, c0_n64_w164, c0_n64_w165, c0_n64_w166, c0_n64_w167, c0_n64_w168, c0_n64_w169, c0_n64_w170, c0_n64_w171, c0_n64_w172, c0_n64_w173, c0_n64_w174, c0_n64_w175, c0_n64_w176, c0_n64_w177, c0_n64_w178, c0_n64_w179, c0_n64_w180, c0_n64_w181, c0_n64_w182, c0_n64_w183, c0_n64_w184, c0_n64_w185, c0_n64_w186, c0_n64_w187, c0_n64_w188, c0_n64_w189, c0_n64_w190, c0_n64_w191, c0_n64_w192, c0_n64_w193, c0_n64_w194, c0_n64_w195, c0_n64_w196, c0_n64_w197, c0_n64_w198, c0_n64_w199, c0_n64_w200, c0_n65_w1, c0_n65_w2, c0_n65_w3, c0_n65_w4, c0_n65_w5, c0_n65_w6, c0_n65_w7, c0_n65_w8, c0_n65_w9, c0_n65_w10, c0_n65_w11, c0_n65_w12, c0_n65_w13, c0_n65_w14, c0_n65_w15, c0_n65_w16, c0_n65_w17, c0_n65_w18, c0_n65_w19, c0_n65_w20, c0_n65_w21, c0_n65_w22, c0_n65_w23, c0_n65_w24, c0_n65_w25, c0_n65_w26, c0_n65_w27, c0_n65_w28, c0_n65_w29, c0_n65_w30, c0_n65_w31, c0_n65_w32, c0_n65_w33, c0_n65_w34, c0_n65_w35, c0_n65_w36, c0_n65_w37, c0_n65_w38, c0_n65_w39, c0_n65_w40, c0_n65_w41, c0_n65_w42, c0_n65_w43, c0_n65_w44, c0_n65_w45, c0_n65_w46, c0_n65_w47, c0_n65_w48, c0_n65_w49, c0_n65_w50, c0_n65_w51, c0_n65_w52, c0_n65_w53, c0_n65_w54, c0_n65_w55, c0_n65_w56, c0_n65_w57, c0_n65_w58, c0_n65_w59, c0_n65_w60, c0_n65_w61, c0_n65_w62, c0_n65_w63, c0_n65_w64, c0_n65_w65, c0_n65_w66, c0_n65_w67, c0_n65_w68, c0_n65_w69, c0_n65_w70, c0_n65_w71, c0_n65_w72, c0_n65_w73, c0_n65_w74, c0_n65_w75, c0_n65_w76, c0_n65_w77, c0_n65_w78, c0_n65_w79, c0_n65_w80, c0_n65_w81, c0_n65_w82, c0_n65_w83, c0_n65_w84, c0_n65_w85, c0_n65_w86, c0_n65_w87, c0_n65_w88, c0_n65_w89, c0_n65_w90, c0_n65_w91, c0_n65_w92, c0_n65_w93, c0_n65_w94, c0_n65_w95, c0_n65_w96, c0_n65_w97, c0_n65_w98, c0_n65_w99, c0_n65_w100, c0_n65_w101, c0_n65_w102, c0_n65_w103, c0_n65_w104, c0_n65_w105, c0_n65_w106, c0_n65_w107, c0_n65_w108, c0_n65_w109, c0_n65_w110, c0_n65_w111, c0_n65_w112, c0_n65_w113, c0_n65_w114, c0_n65_w115, c0_n65_w116, c0_n65_w117, c0_n65_w118, c0_n65_w119, c0_n65_w120, c0_n65_w121, c0_n65_w122, c0_n65_w123, c0_n65_w124, c0_n65_w125, c0_n65_w126, c0_n65_w127, c0_n65_w128, c0_n65_w129, c0_n65_w130, c0_n65_w131, c0_n65_w132, c0_n65_w133, c0_n65_w134, c0_n65_w135, c0_n65_w136, c0_n65_w137, c0_n65_w138, c0_n65_w139, c0_n65_w140, c0_n65_w141, c0_n65_w142, c0_n65_w143, c0_n65_w144, c0_n65_w145, c0_n65_w146, c0_n65_w147, c0_n65_w148, c0_n65_w149, c0_n65_w150, c0_n65_w151, c0_n65_w152, c0_n65_w153, c0_n65_w154, c0_n65_w155, c0_n65_w156, c0_n65_w157, c0_n65_w158, c0_n65_w159, c0_n65_w160, c0_n65_w161, c0_n65_w162, c0_n65_w163, c0_n65_w164, c0_n65_w165, c0_n65_w166, c0_n65_w167, c0_n65_w168, c0_n65_w169, c0_n65_w170, c0_n65_w171, c0_n65_w172, c0_n65_w173, c0_n65_w174, c0_n65_w175, c0_n65_w176, c0_n65_w177, c0_n65_w178, c0_n65_w179, c0_n65_w180, c0_n65_w181, c0_n65_w182, c0_n65_w183, c0_n65_w184, c0_n65_w185, c0_n65_w186, c0_n65_w187, c0_n65_w188, c0_n65_w189, c0_n65_w190, c0_n65_w191, c0_n65_w192, c0_n65_w193, c0_n65_w194, c0_n65_w195, c0_n65_w196, c0_n65_w197, c0_n65_w198, c0_n65_w199, c0_n65_w200, c0_n66_w1, c0_n66_w2, c0_n66_w3, c0_n66_w4, c0_n66_w5, c0_n66_w6, c0_n66_w7, c0_n66_w8, c0_n66_w9, c0_n66_w10, c0_n66_w11, c0_n66_w12, c0_n66_w13, c0_n66_w14, c0_n66_w15, c0_n66_w16, c0_n66_w17, c0_n66_w18, c0_n66_w19, c0_n66_w20, c0_n66_w21, c0_n66_w22, c0_n66_w23, c0_n66_w24, c0_n66_w25, c0_n66_w26, c0_n66_w27, c0_n66_w28, c0_n66_w29, c0_n66_w30, c0_n66_w31, c0_n66_w32, c0_n66_w33, c0_n66_w34, c0_n66_w35, c0_n66_w36, c0_n66_w37, c0_n66_w38, c0_n66_w39, c0_n66_w40, c0_n66_w41, c0_n66_w42, c0_n66_w43, c0_n66_w44, c0_n66_w45, c0_n66_w46, c0_n66_w47, c0_n66_w48, c0_n66_w49, c0_n66_w50, c0_n66_w51, c0_n66_w52, c0_n66_w53, c0_n66_w54, c0_n66_w55, c0_n66_w56, c0_n66_w57, c0_n66_w58, c0_n66_w59, c0_n66_w60, c0_n66_w61, c0_n66_w62, c0_n66_w63, c0_n66_w64, c0_n66_w65, c0_n66_w66, c0_n66_w67, c0_n66_w68, c0_n66_w69, c0_n66_w70, c0_n66_w71, c0_n66_w72, c0_n66_w73, c0_n66_w74, c0_n66_w75, c0_n66_w76, c0_n66_w77, c0_n66_w78, c0_n66_w79, c0_n66_w80, c0_n66_w81, c0_n66_w82, c0_n66_w83, c0_n66_w84, c0_n66_w85, c0_n66_w86, c0_n66_w87, c0_n66_w88, c0_n66_w89, c0_n66_w90, c0_n66_w91, c0_n66_w92, c0_n66_w93, c0_n66_w94, c0_n66_w95, c0_n66_w96, c0_n66_w97, c0_n66_w98, c0_n66_w99, c0_n66_w100, c0_n66_w101, c0_n66_w102, c0_n66_w103, c0_n66_w104, c0_n66_w105, c0_n66_w106, c0_n66_w107, c0_n66_w108, c0_n66_w109, c0_n66_w110, c0_n66_w111, c0_n66_w112, c0_n66_w113, c0_n66_w114, c0_n66_w115, c0_n66_w116, c0_n66_w117, c0_n66_w118, c0_n66_w119, c0_n66_w120, c0_n66_w121, c0_n66_w122, c0_n66_w123, c0_n66_w124, c0_n66_w125, c0_n66_w126, c0_n66_w127, c0_n66_w128, c0_n66_w129, c0_n66_w130, c0_n66_w131, c0_n66_w132, c0_n66_w133, c0_n66_w134, c0_n66_w135, c0_n66_w136, c0_n66_w137, c0_n66_w138, c0_n66_w139, c0_n66_w140, c0_n66_w141, c0_n66_w142, c0_n66_w143, c0_n66_w144, c0_n66_w145, c0_n66_w146, c0_n66_w147, c0_n66_w148, c0_n66_w149, c0_n66_w150, c0_n66_w151, c0_n66_w152, c0_n66_w153, c0_n66_w154, c0_n66_w155, c0_n66_w156, c0_n66_w157, c0_n66_w158, c0_n66_w159, c0_n66_w160, c0_n66_w161, c0_n66_w162, c0_n66_w163, c0_n66_w164, c0_n66_w165, c0_n66_w166, c0_n66_w167, c0_n66_w168, c0_n66_w169, c0_n66_w170, c0_n66_w171, c0_n66_w172, c0_n66_w173, c0_n66_w174, c0_n66_w175, c0_n66_w176, c0_n66_w177, c0_n66_w178, c0_n66_w179, c0_n66_w180, c0_n66_w181, c0_n66_w182, c0_n66_w183, c0_n66_w184, c0_n66_w185, c0_n66_w186, c0_n66_w187, c0_n66_w188, c0_n66_w189, c0_n66_w190, c0_n66_w191, c0_n66_w192, c0_n66_w193, c0_n66_w194, c0_n66_w195, c0_n66_w196, c0_n66_w197, c0_n66_w198, c0_n66_w199, c0_n66_w200, c0_n67_w1, c0_n67_w2, c0_n67_w3, c0_n67_w4, c0_n67_w5, c0_n67_w6, c0_n67_w7, c0_n67_w8, c0_n67_w9, c0_n67_w10, c0_n67_w11, c0_n67_w12, c0_n67_w13, c0_n67_w14, c0_n67_w15, c0_n67_w16, c0_n67_w17, c0_n67_w18, c0_n67_w19, c0_n67_w20, c0_n67_w21, c0_n67_w22, c0_n67_w23, c0_n67_w24, c0_n67_w25, c0_n67_w26, c0_n67_w27, c0_n67_w28, c0_n67_w29, c0_n67_w30, c0_n67_w31, c0_n67_w32, c0_n67_w33, c0_n67_w34, c0_n67_w35, c0_n67_w36, c0_n67_w37, c0_n67_w38, c0_n67_w39, c0_n67_w40, c0_n67_w41, c0_n67_w42, c0_n67_w43, c0_n67_w44, c0_n67_w45, c0_n67_w46, c0_n67_w47, c0_n67_w48, c0_n67_w49, c0_n67_w50, c0_n67_w51, c0_n67_w52, c0_n67_w53, c0_n67_w54, c0_n67_w55, c0_n67_w56, c0_n67_w57, c0_n67_w58, c0_n67_w59, c0_n67_w60, c0_n67_w61, c0_n67_w62, c0_n67_w63, c0_n67_w64, c0_n67_w65, c0_n67_w66, c0_n67_w67, c0_n67_w68, c0_n67_w69, c0_n67_w70, c0_n67_w71, c0_n67_w72, c0_n67_w73, c0_n67_w74, c0_n67_w75, c0_n67_w76, c0_n67_w77, c0_n67_w78, c0_n67_w79, c0_n67_w80, c0_n67_w81, c0_n67_w82, c0_n67_w83, c0_n67_w84, c0_n67_w85, c0_n67_w86, c0_n67_w87, c0_n67_w88, c0_n67_w89, c0_n67_w90, c0_n67_w91, c0_n67_w92, c0_n67_w93, c0_n67_w94, c0_n67_w95, c0_n67_w96, c0_n67_w97, c0_n67_w98, c0_n67_w99, c0_n67_w100, c0_n67_w101, c0_n67_w102, c0_n67_w103, c0_n67_w104, c0_n67_w105, c0_n67_w106, c0_n67_w107, c0_n67_w108, c0_n67_w109, c0_n67_w110, c0_n67_w111, c0_n67_w112, c0_n67_w113, c0_n67_w114, c0_n67_w115, c0_n67_w116, c0_n67_w117, c0_n67_w118, c0_n67_w119, c0_n67_w120, c0_n67_w121, c0_n67_w122, c0_n67_w123, c0_n67_w124, c0_n67_w125, c0_n67_w126, c0_n67_w127, c0_n67_w128, c0_n67_w129, c0_n67_w130, c0_n67_w131, c0_n67_w132, c0_n67_w133, c0_n67_w134, c0_n67_w135, c0_n67_w136, c0_n67_w137, c0_n67_w138, c0_n67_w139, c0_n67_w140, c0_n67_w141, c0_n67_w142, c0_n67_w143, c0_n67_w144, c0_n67_w145, c0_n67_w146, c0_n67_w147, c0_n67_w148, c0_n67_w149, c0_n67_w150, c0_n67_w151, c0_n67_w152, c0_n67_w153, c0_n67_w154, c0_n67_w155, c0_n67_w156, c0_n67_w157, c0_n67_w158, c0_n67_w159, c0_n67_w160, c0_n67_w161, c0_n67_w162, c0_n67_w163, c0_n67_w164, c0_n67_w165, c0_n67_w166, c0_n67_w167, c0_n67_w168, c0_n67_w169, c0_n67_w170, c0_n67_w171, c0_n67_w172, c0_n67_w173, c0_n67_w174, c0_n67_w175, c0_n67_w176, c0_n67_w177, c0_n67_w178, c0_n67_w179, c0_n67_w180, c0_n67_w181, c0_n67_w182, c0_n67_w183, c0_n67_w184, c0_n67_w185, c0_n67_w186, c0_n67_w187, c0_n67_w188, c0_n67_w189, c0_n67_w190, c0_n67_w191, c0_n67_w192, c0_n67_w193, c0_n67_w194, c0_n67_w195, c0_n67_w196, c0_n67_w197, c0_n67_w198, c0_n67_w199, c0_n67_w200, c0_n68_w1, c0_n68_w2, c0_n68_w3, c0_n68_w4, c0_n68_w5, c0_n68_w6, c0_n68_w7, c0_n68_w8, c0_n68_w9, c0_n68_w10, c0_n68_w11, c0_n68_w12, c0_n68_w13, c0_n68_w14, c0_n68_w15, c0_n68_w16, c0_n68_w17, c0_n68_w18, c0_n68_w19, c0_n68_w20, c0_n68_w21, c0_n68_w22, c0_n68_w23, c0_n68_w24, c0_n68_w25, c0_n68_w26, c0_n68_w27, c0_n68_w28, c0_n68_w29, c0_n68_w30, c0_n68_w31, c0_n68_w32, c0_n68_w33, c0_n68_w34, c0_n68_w35, c0_n68_w36, c0_n68_w37, c0_n68_w38, c0_n68_w39, c0_n68_w40, c0_n68_w41, c0_n68_w42, c0_n68_w43, c0_n68_w44, c0_n68_w45, c0_n68_w46, c0_n68_w47, c0_n68_w48, c0_n68_w49, c0_n68_w50, c0_n68_w51, c0_n68_w52, c0_n68_w53, c0_n68_w54, c0_n68_w55, c0_n68_w56, c0_n68_w57, c0_n68_w58, c0_n68_w59, c0_n68_w60, c0_n68_w61, c0_n68_w62, c0_n68_w63, c0_n68_w64, c0_n68_w65, c0_n68_w66, c0_n68_w67, c0_n68_w68, c0_n68_w69, c0_n68_w70, c0_n68_w71, c0_n68_w72, c0_n68_w73, c0_n68_w74, c0_n68_w75, c0_n68_w76, c0_n68_w77, c0_n68_w78, c0_n68_w79, c0_n68_w80, c0_n68_w81, c0_n68_w82, c0_n68_w83, c0_n68_w84, c0_n68_w85, c0_n68_w86, c0_n68_w87, c0_n68_w88, c0_n68_w89, c0_n68_w90, c0_n68_w91, c0_n68_w92, c0_n68_w93, c0_n68_w94, c0_n68_w95, c0_n68_w96, c0_n68_w97, c0_n68_w98, c0_n68_w99, c0_n68_w100, c0_n68_w101, c0_n68_w102, c0_n68_w103, c0_n68_w104, c0_n68_w105, c0_n68_w106, c0_n68_w107, c0_n68_w108, c0_n68_w109, c0_n68_w110, c0_n68_w111, c0_n68_w112, c0_n68_w113, c0_n68_w114, c0_n68_w115, c0_n68_w116, c0_n68_w117, c0_n68_w118, c0_n68_w119, c0_n68_w120, c0_n68_w121, c0_n68_w122, c0_n68_w123, c0_n68_w124, c0_n68_w125, c0_n68_w126, c0_n68_w127, c0_n68_w128, c0_n68_w129, c0_n68_w130, c0_n68_w131, c0_n68_w132, c0_n68_w133, c0_n68_w134, c0_n68_w135, c0_n68_w136, c0_n68_w137, c0_n68_w138, c0_n68_w139, c0_n68_w140, c0_n68_w141, c0_n68_w142, c0_n68_w143, c0_n68_w144, c0_n68_w145, c0_n68_w146, c0_n68_w147, c0_n68_w148, c0_n68_w149, c0_n68_w150, c0_n68_w151, c0_n68_w152, c0_n68_w153, c0_n68_w154, c0_n68_w155, c0_n68_w156, c0_n68_w157, c0_n68_w158, c0_n68_w159, c0_n68_w160, c0_n68_w161, c0_n68_w162, c0_n68_w163, c0_n68_w164, c0_n68_w165, c0_n68_w166, c0_n68_w167, c0_n68_w168, c0_n68_w169, c0_n68_w170, c0_n68_w171, c0_n68_w172, c0_n68_w173, c0_n68_w174, c0_n68_w175, c0_n68_w176, c0_n68_w177, c0_n68_w178, c0_n68_w179, c0_n68_w180, c0_n68_w181, c0_n68_w182, c0_n68_w183, c0_n68_w184, c0_n68_w185, c0_n68_w186, c0_n68_w187, c0_n68_w188, c0_n68_w189, c0_n68_w190, c0_n68_w191, c0_n68_w192, c0_n68_w193, c0_n68_w194, c0_n68_w195, c0_n68_w196, c0_n68_w197, c0_n68_w198, c0_n68_w199, c0_n68_w200, c0_n69_w1, c0_n69_w2, c0_n69_w3, c0_n69_w4, c0_n69_w5, c0_n69_w6, c0_n69_w7, c0_n69_w8, c0_n69_w9, c0_n69_w10, c0_n69_w11, c0_n69_w12, c0_n69_w13, c0_n69_w14, c0_n69_w15, c0_n69_w16, c0_n69_w17, c0_n69_w18, c0_n69_w19, c0_n69_w20, c0_n69_w21, c0_n69_w22, c0_n69_w23, c0_n69_w24, c0_n69_w25, c0_n69_w26, c0_n69_w27, c0_n69_w28, c0_n69_w29, c0_n69_w30, c0_n69_w31, c0_n69_w32, c0_n69_w33, c0_n69_w34, c0_n69_w35, c0_n69_w36, c0_n69_w37, c0_n69_w38, c0_n69_w39, c0_n69_w40, c0_n69_w41, c0_n69_w42, c0_n69_w43, c0_n69_w44, c0_n69_w45, c0_n69_w46, c0_n69_w47, c0_n69_w48, c0_n69_w49, c0_n69_w50, c0_n69_w51, c0_n69_w52, c0_n69_w53, c0_n69_w54, c0_n69_w55, c0_n69_w56, c0_n69_w57, c0_n69_w58, c0_n69_w59, c0_n69_w60, c0_n69_w61, c0_n69_w62, c0_n69_w63, c0_n69_w64, c0_n69_w65, c0_n69_w66, c0_n69_w67, c0_n69_w68, c0_n69_w69, c0_n69_w70, c0_n69_w71, c0_n69_w72, c0_n69_w73, c0_n69_w74, c0_n69_w75, c0_n69_w76, c0_n69_w77, c0_n69_w78, c0_n69_w79, c0_n69_w80, c0_n69_w81, c0_n69_w82, c0_n69_w83, c0_n69_w84, c0_n69_w85, c0_n69_w86, c0_n69_w87, c0_n69_w88, c0_n69_w89, c0_n69_w90, c0_n69_w91, c0_n69_w92, c0_n69_w93, c0_n69_w94, c0_n69_w95, c0_n69_w96, c0_n69_w97, c0_n69_w98, c0_n69_w99, c0_n69_w100, c0_n69_w101, c0_n69_w102, c0_n69_w103, c0_n69_w104, c0_n69_w105, c0_n69_w106, c0_n69_w107, c0_n69_w108, c0_n69_w109, c0_n69_w110, c0_n69_w111, c0_n69_w112, c0_n69_w113, c0_n69_w114, c0_n69_w115, c0_n69_w116, c0_n69_w117, c0_n69_w118, c0_n69_w119, c0_n69_w120, c0_n69_w121, c0_n69_w122, c0_n69_w123, c0_n69_w124, c0_n69_w125, c0_n69_w126, c0_n69_w127, c0_n69_w128, c0_n69_w129, c0_n69_w130, c0_n69_w131, c0_n69_w132, c0_n69_w133, c0_n69_w134, c0_n69_w135, c0_n69_w136, c0_n69_w137, c0_n69_w138, c0_n69_w139, c0_n69_w140, c0_n69_w141, c0_n69_w142, c0_n69_w143, c0_n69_w144, c0_n69_w145, c0_n69_w146, c0_n69_w147, c0_n69_w148, c0_n69_w149, c0_n69_w150, c0_n69_w151, c0_n69_w152, c0_n69_w153, c0_n69_w154, c0_n69_w155, c0_n69_w156, c0_n69_w157, c0_n69_w158, c0_n69_w159, c0_n69_w160, c0_n69_w161, c0_n69_w162, c0_n69_w163, c0_n69_w164, c0_n69_w165, c0_n69_w166, c0_n69_w167, c0_n69_w168, c0_n69_w169, c0_n69_w170, c0_n69_w171, c0_n69_w172, c0_n69_w173, c0_n69_w174, c0_n69_w175, c0_n69_w176, c0_n69_w177, c0_n69_w178, c0_n69_w179, c0_n69_w180, c0_n69_w181, c0_n69_w182, c0_n69_w183, c0_n69_w184, c0_n69_w185, c0_n69_w186, c0_n69_w187, c0_n69_w188, c0_n69_w189, c0_n69_w190, c0_n69_w191, c0_n69_w192, c0_n69_w193, c0_n69_w194, c0_n69_w195, c0_n69_w196, c0_n69_w197, c0_n69_w198, c0_n69_w199, c0_n69_w200, c0_n70_w1, c0_n70_w2, c0_n70_w3, c0_n70_w4, c0_n70_w5, c0_n70_w6, c0_n70_w7, c0_n70_w8, c0_n70_w9, c0_n70_w10, c0_n70_w11, c0_n70_w12, c0_n70_w13, c0_n70_w14, c0_n70_w15, c0_n70_w16, c0_n70_w17, c0_n70_w18, c0_n70_w19, c0_n70_w20, c0_n70_w21, c0_n70_w22, c0_n70_w23, c0_n70_w24, c0_n70_w25, c0_n70_w26, c0_n70_w27, c0_n70_w28, c0_n70_w29, c0_n70_w30, c0_n70_w31, c0_n70_w32, c0_n70_w33, c0_n70_w34, c0_n70_w35, c0_n70_w36, c0_n70_w37, c0_n70_w38, c0_n70_w39, c0_n70_w40, c0_n70_w41, c0_n70_w42, c0_n70_w43, c0_n70_w44, c0_n70_w45, c0_n70_w46, c0_n70_w47, c0_n70_w48, c0_n70_w49, c0_n70_w50, c0_n70_w51, c0_n70_w52, c0_n70_w53, c0_n70_w54, c0_n70_w55, c0_n70_w56, c0_n70_w57, c0_n70_w58, c0_n70_w59, c0_n70_w60, c0_n70_w61, c0_n70_w62, c0_n70_w63, c0_n70_w64, c0_n70_w65, c0_n70_w66, c0_n70_w67, c0_n70_w68, c0_n70_w69, c0_n70_w70, c0_n70_w71, c0_n70_w72, c0_n70_w73, c0_n70_w74, c0_n70_w75, c0_n70_w76, c0_n70_w77, c0_n70_w78, c0_n70_w79, c0_n70_w80, c0_n70_w81, c0_n70_w82, c0_n70_w83, c0_n70_w84, c0_n70_w85, c0_n70_w86, c0_n70_w87, c0_n70_w88, c0_n70_w89, c0_n70_w90, c0_n70_w91, c0_n70_w92, c0_n70_w93, c0_n70_w94, c0_n70_w95, c0_n70_w96, c0_n70_w97, c0_n70_w98, c0_n70_w99, c0_n70_w100, c0_n70_w101, c0_n70_w102, c0_n70_w103, c0_n70_w104, c0_n70_w105, c0_n70_w106, c0_n70_w107, c0_n70_w108, c0_n70_w109, c0_n70_w110, c0_n70_w111, c0_n70_w112, c0_n70_w113, c0_n70_w114, c0_n70_w115, c0_n70_w116, c0_n70_w117, c0_n70_w118, c0_n70_w119, c0_n70_w120, c0_n70_w121, c0_n70_w122, c0_n70_w123, c0_n70_w124, c0_n70_w125, c0_n70_w126, c0_n70_w127, c0_n70_w128, c0_n70_w129, c0_n70_w130, c0_n70_w131, c0_n70_w132, c0_n70_w133, c0_n70_w134, c0_n70_w135, c0_n70_w136, c0_n70_w137, c0_n70_w138, c0_n70_w139, c0_n70_w140, c0_n70_w141, c0_n70_w142, c0_n70_w143, c0_n70_w144, c0_n70_w145, c0_n70_w146, c0_n70_w147, c0_n70_w148, c0_n70_w149, c0_n70_w150, c0_n70_w151, c0_n70_w152, c0_n70_w153, c0_n70_w154, c0_n70_w155, c0_n70_w156, c0_n70_w157, c0_n70_w158, c0_n70_w159, c0_n70_w160, c0_n70_w161, c0_n70_w162, c0_n70_w163, c0_n70_w164, c0_n70_w165, c0_n70_w166, c0_n70_w167, c0_n70_w168, c0_n70_w169, c0_n70_w170, c0_n70_w171, c0_n70_w172, c0_n70_w173, c0_n70_w174, c0_n70_w175, c0_n70_w176, c0_n70_w177, c0_n70_w178, c0_n70_w179, c0_n70_w180, c0_n70_w181, c0_n70_w182, c0_n70_w183, c0_n70_w184, c0_n70_w185, c0_n70_w186, c0_n70_w187, c0_n70_w188, c0_n70_w189, c0_n70_w190, c0_n70_w191, c0_n70_w192, c0_n70_w193, c0_n70_w194, c0_n70_w195, c0_n70_w196, c0_n70_w197, c0_n70_w198, c0_n70_w199, c0_n70_w200, c0_n71_w1, c0_n71_w2, c0_n71_w3, c0_n71_w4, c0_n71_w5, c0_n71_w6, c0_n71_w7, c0_n71_w8, c0_n71_w9, c0_n71_w10, c0_n71_w11, c0_n71_w12, c0_n71_w13, c0_n71_w14, c0_n71_w15, c0_n71_w16, c0_n71_w17, c0_n71_w18, c0_n71_w19, c0_n71_w20, c0_n71_w21, c0_n71_w22, c0_n71_w23, c0_n71_w24, c0_n71_w25, c0_n71_w26, c0_n71_w27, c0_n71_w28, c0_n71_w29, c0_n71_w30, c0_n71_w31, c0_n71_w32, c0_n71_w33, c0_n71_w34, c0_n71_w35, c0_n71_w36, c0_n71_w37, c0_n71_w38, c0_n71_w39, c0_n71_w40, c0_n71_w41, c0_n71_w42, c0_n71_w43, c0_n71_w44, c0_n71_w45, c0_n71_w46, c0_n71_w47, c0_n71_w48, c0_n71_w49, c0_n71_w50, c0_n71_w51, c0_n71_w52, c0_n71_w53, c0_n71_w54, c0_n71_w55, c0_n71_w56, c0_n71_w57, c0_n71_w58, c0_n71_w59, c0_n71_w60, c0_n71_w61, c0_n71_w62, c0_n71_w63, c0_n71_w64, c0_n71_w65, c0_n71_w66, c0_n71_w67, c0_n71_w68, c0_n71_w69, c0_n71_w70, c0_n71_w71, c0_n71_w72, c0_n71_w73, c0_n71_w74, c0_n71_w75, c0_n71_w76, c0_n71_w77, c0_n71_w78, c0_n71_w79, c0_n71_w80, c0_n71_w81, c0_n71_w82, c0_n71_w83, c0_n71_w84, c0_n71_w85, c0_n71_w86, c0_n71_w87, c0_n71_w88, c0_n71_w89, c0_n71_w90, c0_n71_w91, c0_n71_w92, c0_n71_w93, c0_n71_w94, c0_n71_w95, c0_n71_w96, c0_n71_w97, c0_n71_w98, c0_n71_w99, c0_n71_w100, c0_n71_w101, c0_n71_w102, c0_n71_w103, c0_n71_w104, c0_n71_w105, c0_n71_w106, c0_n71_w107, c0_n71_w108, c0_n71_w109, c0_n71_w110, c0_n71_w111, c0_n71_w112, c0_n71_w113, c0_n71_w114, c0_n71_w115, c0_n71_w116, c0_n71_w117, c0_n71_w118, c0_n71_w119, c0_n71_w120, c0_n71_w121, c0_n71_w122, c0_n71_w123, c0_n71_w124, c0_n71_w125, c0_n71_w126, c0_n71_w127, c0_n71_w128, c0_n71_w129, c0_n71_w130, c0_n71_w131, c0_n71_w132, c0_n71_w133, c0_n71_w134, c0_n71_w135, c0_n71_w136, c0_n71_w137, c0_n71_w138, c0_n71_w139, c0_n71_w140, c0_n71_w141, c0_n71_w142, c0_n71_w143, c0_n71_w144, c0_n71_w145, c0_n71_w146, c0_n71_w147, c0_n71_w148, c0_n71_w149, c0_n71_w150, c0_n71_w151, c0_n71_w152, c0_n71_w153, c0_n71_w154, c0_n71_w155, c0_n71_w156, c0_n71_w157, c0_n71_w158, c0_n71_w159, c0_n71_w160, c0_n71_w161, c0_n71_w162, c0_n71_w163, c0_n71_w164, c0_n71_w165, c0_n71_w166, c0_n71_w167, c0_n71_w168, c0_n71_w169, c0_n71_w170, c0_n71_w171, c0_n71_w172, c0_n71_w173, c0_n71_w174, c0_n71_w175, c0_n71_w176, c0_n71_w177, c0_n71_w178, c0_n71_w179, c0_n71_w180, c0_n71_w181, c0_n71_w182, c0_n71_w183, c0_n71_w184, c0_n71_w185, c0_n71_w186, c0_n71_w187, c0_n71_w188, c0_n71_w189, c0_n71_w190, c0_n71_w191, c0_n71_w192, c0_n71_w193, c0_n71_w194, c0_n71_w195, c0_n71_w196, c0_n71_w197, c0_n71_w198, c0_n71_w199, c0_n71_w200, c0_n72_w1, c0_n72_w2, c0_n72_w3, c0_n72_w4, c0_n72_w5, c0_n72_w6, c0_n72_w7, c0_n72_w8, c0_n72_w9, c0_n72_w10, c0_n72_w11, c0_n72_w12, c0_n72_w13, c0_n72_w14, c0_n72_w15, c0_n72_w16, c0_n72_w17, c0_n72_w18, c0_n72_w19, c0_n72_w20, c0_n72_w21, c0_n72_w22, c0_n72_w23, c0_n72_w24, c0_n72_w25, c0_n72_w26, c0_n72_w27, c0_n72_w28, c0_n72_w29, c0_n72_w30, c0_n72_w31, c0_n72_w32, c0_n72_w33, c0_n72_w34, c0_n72_w35, c0_n72_w36, c0_n72_w37, c0_n72_w38, c0_n72_w39, c0_n72_w40, c0_n72_w41, c0_n72_w42, c0_n72_w43, c0_n72_w44, c0_n72_w45, c0_n72_w46, c0_n72_w47, c0_n72_w48, c0_n72_w49, c0_n72_w50, c0_n72_w51, c0_n72_w52, c0_n72_w53, c0_n72_w54, c0_n72_w55, c0_n72_w56, c0_n72_w57, c0_n72_w58, c0_n72_w59, c0_n72_w60, c0_n72_w61, c0_n72_w62, c0_n72_w63, c0_n72_w64, c0_n72_w65, c0_n72_w66, c0_n72_w67, c0_n72_w68, c0_n72_w69, c0_n72_w70, c0_n72_w71, c0_n72_w72, c0_n72_w73, c0_n72_w74, c0_n72_w75, c0_n72_w76, c0_n72_w77, c0_n72_w78, c0_n72_w79, c0_n72_w80, c0_n72_w81, c0_n72_w82, c0_n72_w83, c0_n72_w84, c0_n72_w85, c0_n72_w86, c0_n72_w87, c0_n72_w88, c0_n72_w89, c0_n72_w90, c0_n72_w91, c0_n72_w92, c0_n72_w93, c0_n72_w94, c0_n72_w95, c0_n72_w96, c0_n72_w97, c0_n72_w98, c0_n72_w99, c0_n72_w100, c0_n72_w101, c0_n72_w102, c0_n72_w103, c0_n72_w104, c0_n72_w105, c0_n72_w106, c0_n72_w107, c0_n72_w108, c0_n72_w109, c0_n72_w110, c0_n72_w111, c0_n72_w112, c0_n72_w113, c0_n72_w114, c0_n72_w115, c0_n72_w116, c0_n72_w117, c0_n72_w118, c0_n72_w119, c0_n72_w120, c0_n72_w121, c0_n72_w122, c0_n72_w123, c0_n72_w124, c0_n72_w125, c0_n72_w126, c0_n72_w127, c0_n72_w128, c0_n72_w129, c0_n72_w130, c0_n72_w131, c0_n72_w132, c0_n72_w133, c0_n72_w134, c0_n72_w135, c0_n72_w136, c0_n72_w137, c0_n72_w138, c0_n72_w139, c0_n72_w140, c0_n72_w141, c0_n72_w142, c0_n72_w143, c0_n72_w144, c0_n72_w145, c0_n72_w146, c0_n72_w147, c0_n72_w148, c0_n72_w149, c0_n72_w150, c0_n72_w151, c0_n72_w152, c0_n72_w153, c0_n72_w154, c0_n72_w155, c0_n72_w156, c0_n72_w157, c0_n72_w158, c0_n72_w159, c0_n72_w160, c0_n72_w161, c0_n72_w162, c0_n72_w163, c0_n72_w164, c0_n72_w165, c0_n72_w166, c0_n72_w167, c0_n72_w168, c0_n72_w169, c0_n72_w170, c0_n72_w171, c0_n72_w172, c0_n72_w173, c0_n72_w174, c0_n72_w175, c0_n72_w176, c0_n72_w177, c0_n72_w178, c0_n72_w179, c0_n72_w180, c0_n72_w181, c0_n72_w182, c0_n72_w183, c0_n72_w184, c0_n72_w185, c0_n72_w186, c0_n72_w187, c0_n72_w188, c0_n72_w189, c0_n72_w190, c0_n72_w191, c0_n72_w192, c0_n72_w193, c0_n72_w194, c0_n72_w195, c0_n72_w196, c0_n72_w197, c0_n72_w198, c0_n72_w199, c0_n72_w200, c0_n73_w1, c0_n73_w2, c0_n73_w3, c0_n73_w4, c0_n73_w5, c0_n73_w6, c0_n73_w7, c0_n73_w8, c0_n73_w9, c0_n73_w10, c0_n73_w11, c0_n73_w12, c0_n73_w13, c0_n73_w14, c0_n73_w15, c0_n73_w16, c0_n73_w17, c0_n73_w18, c0_n73_w19, c0_n73_w20, c0_n73_w21, c0_n73_w22, c0_n73_w23, c0_n73_w24, c0_n73_w25, c0_n73_w26, c0_n73_w27, c0_n73_w28, c0_n73_w29, c0_n73_w30, c0_n73_w31, c0_n73_w32, c0_n73_w33, c0_n73_w34, c0_n73_w35, c0_n73_w36, c0_n73_w37, c0_n73_w38, c0_n73_w39, c0_n73_w40, c0_n73_w41, c0_n73_w42, c0_n73_w43, c0_n73_w44, c0_n73_w45, c0_n73_w46, c0_n73_w47, c0_n73_w48, c0_n73_w49, c0_n73_w50, c0_n73_w51, c0_n73_w52, c0_n73_w53, c0_n73_w54, c0_n73_w55, c0_n73_w56, c0_n73_w57, c0_n73_w58, c0_n73_w59, c0_n73_w60, c0_n73_w61, c0_n73_w62, c0_n73_w63, c0_n73_w64, c0_n73_w65, c0_n73_w66, c0_n73_w67, c0_n73_w68, c0_n73_w69, c0_n73_w70, c0_n73_w71, c0_n73_w72, c0_n73_w73, c0_n73_w74, c0_n73_w75, c0_n73_w76, c0_n73_w77, c0_n73_w78, c0_n73_w79, c0_n73_w80, c0_n73_w81, c0_n73_w82, c0_n73_w83, c0_n73_w84, c0_n73_w85, c0_n73_w86, c0_n73_w87, c0_n73_w88, c0_n73_w89, c0_n73_w90, c0_n73_w91, c0_n73_w92, c0_n73_w93, c0_n73_w94, c0_n73_w95, c0_n73_w96, c0_n73_w97, c0_n73_w98, c0_n73_w99, c0_n73_w100, c0_n73_w101, c0_n73_w102, c0_n73_w103, c0_n73_w104, c0_n73_w105, c0_n73_w106, c0_n73_w107, c0_n73_w108, c0_n73_w109, c0_n73_w110, c0_n73_w111, c0_n73_w112, c0_n73_w113, c0_n73_w114, c0_n73_w115, c0_n73_w116, c0_n73_w117, c0_n73_w118, c0_n73_w119, c0_n73_w120, c0_n73_w121, c0_n73_w122, c0_n73_w123, c0_n73_w124, c0_n73_w125, c0_n73_w126, c0_n73_w127, c0_n73_w128, c0_n73_w129, c0_n73_w130, c0_n73_w131, c0_n73_w132, c0_n73_w133, c0_n73_w134, c0_n73_w135, c0_n73_w136, c0_n73_w137, c0_n73_w138, c0_n73_w139, c0_n73_w140, c0_n73_w141, c0_n73_w142, c0_n73_w143, c0_n73_w144, c0_n73_w145, c0_n73_w146, c0_n73_w147, c0_n73_w148, c0_n73_w149, c0_n73_w150, c0_n73_w151, c0_n73_w152, c0_n73_w153, c0_n73_w154, c0_n73_w155, c0_n73_w156, c0_n73_w157, c0_n73_w158, c0_n73_w159, c0_n73_w160, c0_n73_w161, c0_n73_w162, c0_n73_w163, c0_n73_w164, c0_n73_w165, c0_n73_w166, c0_n73_w167, c0_n73_w168, c0_n73_w169, c0_n73_w170, c0_n73_w171, c0_n73_w172, c0_n73_w173, c0_n73_w174, c0_n73_w175, c0_n73_w176, c0_n73_w177, c0_n73_w178, c0_n73_w179, c0_n73_w180, c0_n73_w181, c0_n73_w182, c0_n73_w183, c0_n73_w184, c0_n73_w185, c0_n73_w186, c0_n73_w187, c0_n73_w188, c0_n73_w189, c0_n73_w190, c0_n73_w191, c0_n73_w192, c0_n73_w193, c0_n73_w194, c0_n73_w195, c0_n73_w196, c0_n73_w197, c0_n73_w198, c0_n73_w199, c0_n73_w200, c0_n74_w1, c0_n74_w2, c0_n74_w3, c0_n74_w4, c0_n74_w5, c0_n74_w6, c0_n74_w7, c0_n74_w8, c0_n74_w9, c0_n74_w10, c0_n74_w11, c0_n74_w12, c0_n74_w13, c0_n74_w14, c0_n74_w15, c0_n74_w16, c0_n74_w17, c0_n74_w18, c0_n74_w19, c0_n74_w20, c0_n74_w21, c0_n74_w22, c0_n74_w23, c0_n74_w24, c0_n74_w25, c0_n74_w26, c0_n74_w27, c0_n74_w28, c0_n74_w29, c0_n74_w30, c0_n74_w31, c0_n74_w32, c0_n74_w33, c0_n74_w34, c0_n74_w35, c0_n74_w36, c0_n74_w37, c0_n74_w38, c0_n74_w39, c0_n74_w40, c0_n74_w41, c0_n74_w42, c0_n74_w43, c0_n74_w44, c0_n74_w45, c0_n74_w46, c0_n74_w47, c0_n74_w48, c0_n74_w49, c0_n74_w50, c0_n74_w51, c0_n74_w52, c0_n74_w53, c0_n74_w54, c0_n74_w55, c0_n74_w56, c0_n74_w57, c0_n74_w58, c0_n74_w59, c0_n74_w60, c0_n74_w61, c0_n74_w62, c0_n74_w63, c0_n74_w64, c0_n74_w65, c0_n74_w66, c0_n74_w67, c0_n74_w68, c0_n74_w69, c0_n74_w70, c0_n74_w71, c0_n74_w72, c0_n74_w73, c0_n74_w74, c0_n74_w75, c0_n74_w76, c0_n74_w77, c0_n74_w78, c0_n74_w79, c0_n74_w80, c0_n74_w81, c0_n74_w82, c0_n74_w83, c0_n74_w84, c0_n74_w85, c0_n74_w86, c0_n74_w87, c0_n74_w88, c0_n74_w89, c0_n74_w90, c0_n74_w91, c0_n74_w92, c0_n74_w93, c0_n74_w94, c0_n74_w95, c0_n74_w96, c0_n74_w97, c0_n74_w98, c0_n74_w99, c0_n74_w100, c0_n74_w101, c0_n74_w102, c0_n74_w103, c0_n74_w104, c0_n74_w105, c0_n74_w106, c0_n74_w107, c0_n74_w108, c0_n74_w109, c0_n74_w110, c0_n74_w111, c0_n74_w112, c0_n74_w113, c0_n74_w114, c0_n74_w115, c0_n74_w116, c0_n74_w117, c0_n74_w118, c0_n74_w119, c0_n74_w120, c0_n74_w121, c0_n74_w122, c0_n74_w123, c0_n74_w124, c0_n74_w125, c0_n74_w126, c0_n74_w127, c0_n74_w128, c0_n74_w129, c0_n74_w130, c0_n74_w131, c0_n74_w132, c0_n74_w133, c0_n74_w134, c0_n74_w135, c0_n74_w136, c0_n74_w137, c0_n74_w138, c0_n74_w139, c0_n74_w140, c0_n74_w141, c0_n74_w142, c0_n74_w143, c0_n74_w144, c0_n74_w145, c0_n74_w146, c0_n74_w147, c0_n74_w148, c0_n74_w149, c0_n74_w150, c0_n74_w151, c0_n74_w152, c0_n74_w153, c0_n74_w154, c0_n74_w155, c0_n74_w156, c0_n74_w157, c0_n74_w158, c0_n74_w159, c0_n74_w160, c0_n74_w161, c0_n74_w162, c0_n74_w163, c0_n74_w164, c0_n74_w165, c0_n74_w166, c0_n74_w167, c0_n74_w168, c0_n74_w169, c0_n74_w170, c0_n74_w171, c0_n74_w172, c0_n74_w173, c0_n74_w174, c0_n74_w175, c0_n74_w176, c0_n74_w177, c0_n74_w178, c0_n74_w179, c0_n74_w180, c0_n74_w181, c0_n74_w182, c0_n74_w183, c0_n74_w184, c0_n74_w185, c0_n74_w186, c0_n74_w187, c0_n74_w188, c0_n74_w189, c0_n74_w190, c0_n74_w191, c0_n74_w192, c0_n74_w193, c0_n74_w194, c0_n74_w195, c0_n74_w196, c0_n74_w197, c0_n74_w198, c0_n74_w199, c0_n74_w200, c0_n75_w1, c0_n75_w2, c0_n75_w3, c0_n75_w4, c0_n75_w5, c0_n75_w6, c0_n75_w7, c0_n75_w8, c0_n75_w9, c0_n75_w10, c0_n75_w11, c0_n75_w12, c0_n75_w13, c0_n75_w14, c0_n75_w15, c0_n75_w16, c0_n75_w17, c0_n75_w18, c0_n75_w19, c0_n75_w20, c0_n75_w21, c0_n75_w22, c0_n75_w23, c0_n75_w24, c0_n75_w25, c0_n75_w26, c0_n75_w27, c0_n75_w28, c0_n75_w29, c0_n75_w30, c0_n75_w31, c0_n75_w32, c0_n75_w33, c0_n75_w34, c0_n75_w35, c0_n75_w36, c0_n75_w37, c0_n75_w38, c0_n75_w39, c0_n75_w40, c0_n75_w41, c0_n75_w42, c0_n75_w43, c0_n75_w44, c0_n75_w45, c0_n75_w46, c0_n75_w47, c0_n75_w48, c0_n75_w49, c0_n75_w50, c0_n75_w51, c0_n75_w52, c0_n75_w53, c0_n75_w54, c0_n75_w55, c0_n75_w56, c0_n75_w57, c0_n75_w58, c0_n75_w59, c0_n75_w60, c0_n75_w61, c0_n75_w62, c0_n75_w63, c0_n75_w64, c0_n75_w65, c0_n75_w66, c0_n75_w67, c0_n75_w68, c0_n75_w69, c0_n75_w70, c0_n75_w71, c0_n75_w72, c0_n75_w73, c0_n75_w74, c0_n75_w75, c0_n75_w76, c0_n75_w77, c0_n75_w78, c0_n75_w79, c0_n75_w80, c0_n75_w81, c0_n75_w82, c0_n75_w83, c0_n75_w84, c0_n75_w85, c0_n75_w86, c0_n75_w87, c0_n75_w88, c0_n75_w89, c0_n75_w90, c0_n75_w91, c0_n75_w92, c0_n75_w93, c0_n75_w94, c0_n75_w95, c0_n75_w96, c0_n75_w97, c0_n75_w98, c0_n75_w99, c0_n75_w100, c0_n75_w101, c0_n75_w102, c0_n75_w103, c0_n75_w104, c0_n75_w105, c0_n75_w106, c0_n75_w107, c0_n75_w108, c0_n75_w109, c0_n75_w110, c0_n75_w111, c0_n75_w112, c0_n75_w113, c0_n75_w114, c0_n75_w115, c0_n75_w116, c0_n75_w117, c0_n75_w118, c0_n75_w119, c0_n75_w120, c0_n75_w121, c0_n75_w122, c0_n75_w123, c0_n75_w124, c0_n75_w125, c0_n75_w126, c0_n75_w127, c0_n75_w128, c0_n75_w129, c0_n75_w130, c0_n75_w131, c0_n75_w132, c0_n75_w133, c0_n75_w134, c0_n75_w135, c0_n75_w136, c0_n75_w137, c0_n75_w138, c0_n75_w139, c0_n75_w140, c0_n75_w141, c0_n75_w142, c0_n75_w143, c0_n75_w144, c0_n75_w145, c0_n75_w146, c0_n75_w147, c0_n75_w148, c0_n75_w149, c0_n75_w150, c0_n75_w151, c0_n75_w152, c0_n75_w153, c0_n75_w154, c0_n75_w155, c0_n75_w156, c0_n75_w157, c0_n75_w158, c0_n75_w159, c0_n75_w160, c0_n75_w161, c0_n75_w162, c0_n75_w163, c0_n75_w164, c0_n75_w165, c0_n75_w166, c0_n75_w167, c0_n75_w168, c0_n75_w169, c0_n75_w170, c0_n75_w171, c0_n75_w172, c0_n75_w173, c0_n75_w174, c0_n75_w175, c0_n75_w176, c0_n75_w177, c0_n75_w178, c0_n75_w179, c0_n75_w180, c0_n75_w181, c0_n75_w182, c0_n75_w183, c0_n75_w184, c0_n75_w185, c0_n75_w186, c0_n75_w187, c0_n75_w188, c0_n75_w189, c0_n75_w190, c0_n75_w191, c0_n75_w192, c0_n75_w193, c0_n75_w194, c0_n75_w195, c0_n75_w196, c0_n75_w197, c0_n75_w198, c0_n75_w199, c0_n75_w200, c0_n76_w1, c0_n76_w2, c0_n76_w3, c0_n76_w4, c0_n76_w5, c0_n76_w6, c0_n76_w7, c0_n76_w8, c0_n76_w9, c0_n76_w10, c0_n76_w11, c0_n76_w12, c0_n76_w13, c0_n76_w14, c0_n76_w15, c0_n76_w16, c0_n76_w17, c0_n76_w18, c0_n76_w19, c0_n76_w20, c0_n76_w21, c0_n76_w22, c0_n76_w23, c0_n76_w24, c0_n76_w25, c0_n76_w26, c0_n76_w27, c0_n76_w28, c0_n76_w29, c0_n76_w30, c0_n76_w31, c0_n76_w32, c0_n76_w33, c0_n76_w34, c0_n76_w35, c0_n76_w36, c0_n76_w37, c0_n76_w38, c0_n76_w39, c0_n76_w40, c0_n76_w41, c0_n76_w42, c0_n76_w43, c0_n76_w44, c0_n76_w45, c0_n76_w46, c0_n76_w47, c0_n76_w48, c0_n76_w49, c0_n76_w50, c0_n76_w51, c0_n76_w52, c0_n76_w53, c0_n76_w54, c0_n76_w55, c0_n76_w56, c0_n76_w57, c0_n76_w58, c0_n76_w59, c0_n76_w60, c0_n76_w61, c0_n76_w62, c0_n76_w63, c0_n76_w64, c0_n76_w65, c0_n76_w66, c0_n76_w67, c0_n76_w68, c0_n76_w69, c0_n76_w70, c0_n76_w71, c0_n76_w72, c0_n76_w73, c0_n76_w74, c0_n76_w75, c0_n76_w76, c0_n76_w77, c0_n76_w78, c0_n76_w79, c0_n76_w80, c0_n76_w81, c0_n76_w82, c0_n76_w83, c0_n76_w84, c0_n76_w85, c0_n76_w86, c0_n76_w87, c0_n76_w88, c0_n76_w89, c0_n76_w90, c0_n76_w91, c0_n76_w92, c0_n76_w93, c0_n76_w94, c0_n76_w95, c0_n76_w96, c0_n76_w97, c0_n76_w98, c0_n76_w99, c0_n76_w100, c0_n76_w101, c0_n76_w102, c0_n76_w103, c0_n76_w104, c0_n76_w105, c0_n76_w106, c0_n76_w107, c0_n76_w108, c0_n76_w109, c0_n76_w110, c0_n76_w111, c0_n76_w112, c0_n76_w113, c0_n76_w114, c0_n76_w115, c0_n76_w116, c0_n76_w117, c0_n76_w118, c0_n76_w119, c0_n76_w120, c0_n76_w121, c0_n76_w122, c0_n76_w123, c0_n76_w124, c0_n76_w125, c0_n76_w126, c0_n76_w127, c0_n76_w128, c0_n76_w129, c0_n76_w130, c0_n76_w131, c0_n76_w132, c0_n76_w133, c0_n76_w134, c0_n76_w135, c0_n76_w136, c0_n76_w137, c0_n76_w138, c0_n76_w139, c0_n76_w140, c0_n76_w141, c0_n76_w142, c0_n76_w143, c0_n76_w144, c0_n76_w145, c0_n76_w146, c0_n76_w147, c0_n76_w148, c0_n76_w149, c0_n76_w150, c0_n76_w151, c0_n76_w152, c0_n76_w153, c0_n76_w154, c0_n76_w155, c0_n76_w156, c0_n76_w157, c0_n76_w158, c0_n76_w159, c0_n76_w160, c0_n76_w161, c0_n76_w162, c0_n76_w163, c0_n76_w164, c0_n76_w165, c0_n76_w166, c0_n76_w167, c0_n76_w168, c0_n76_w169, c0_n76_w170, c0_n76_w171, c0_n76_w172, c0_n76_w173, c0_n76_w174, c0_n76_w175, c0_n76_w176, c0_n76_w177, c0_n76_w178, c0_n76_w179, c0_n76_w180, c0_n76_w181, c0_n76_w182, c0_n76_w183, c0_n76_w184, c0_n76_w185, c0_n76_w186, c0_n76_w187, c0_n76_w188, c0_n76_w189, c0_n76_w190, c0_n76_w191, c0_n76_w192, c0_n76_w193, c0_n76_w194, c0_n76_w195, c0_n76_w196, c0_n76_w197, c0_n76_w198, c0_n76_w199, c0_n76_w200, c0_n77_w1, c0_n77_w2, c0_n77_w3, c0_n77_w4, c0_n77_w5, c0_n77_w6, c0_n77_w7, c0_n77_w8, c0_n77_w9, c0_n77_w10, c0_n77_w11, c0_n77_w12, c0_n77_w13, c0_n77_w14, c0_n77_w15, c0_n77_w16, c0_n77_w17, c0_n77_w18, c0_n77_w19, c0_n77_w20, c0_n77_w21, c0_n77_w22, c0_n77_w23, c0_n77_w24, c0_n77_w25, c0_n77_w26, c0_n77_w27, c0_n77_w28, c0_n77_w29, c0_n77_w30, c0_n77_w31, c0_n77_w32, c0_n77_w33, c0_n77_w34, c0_n77_w35, c0_n77_w36, c0_n77_w37, c0_n77_w38, c0_n77_w39, c0_n77_w40, c0_n77_w41, c0_n77_w42, c0_n77_w43, c0_n77_w44, c0_n77_w45, c0_n77_w46, c0_n77_w47, c0_n77_w48, c0_n77_w49, c0_n77_w50, c0_n77_w51, c0_n77_w52, c0_n77_w53, c0_n77_w54, c0_n77_w55, c0_n77_w56, c0_n77_w57, c0_n77_w58, c0_n77_w59, c0_n77_w60, c0_n77_w61, c0_n77_w62, c0_n77_w63, c0_n77_w64, c0_n77_w65, c0_n77_w66, c0_n77_w67, c0_n77_w68, c0_n77_w69, c0_n77_w70, c0_n77_w71, c0_n77_w72, c0_n77_w73, c0_n77_w74, c0_n77_w75, c0_n77_w76, c0_n77_w77, c0_n77_w78, c0_n77_w79, c0_n77_w80, c0_n77_w81, c0_n77_w82, c0_n77_w83, c0_n77_w84, c0_n77_w85, c0_n77_w86, c0_n77_w87, c0_n77_w88, c0_n77_w89, c0_n77_w90, c0_n77_w91, c0_n77_w92, c0_n77_w93, c0_n77_w94, c0_n77_w95, c0_n77_w96, c0_n77_w97, c0_n77_w98, c0_n77_w99, c0_n77_w100, c0_n77_w101, c0_n77_w102, c0_n77_w103, c0_n77_w104, c0_n77_w105, c0_n77_w106, c0_n77_w107, c0_n77_w108, c0_n77_w109, c0_n77_w110, c0_n77_w111, c0_n77_w112, c0_n77_w113, c0_n77_w114, c0_n77_w115, c0_n77_w116, c0_n77_w117, c0_n77_w118, c0_n77_w119, c0_n77_w120, c0_n77_w121, c0_n77_w122, c0_n77_w123, c0_n77_w124, c0_n77_w125, c0_n77_w126, c0_n77_w127, c0_n77_w128, c0_n77_w129, c0_n77_w130, c0_n77_w131, c0_n77_w132, c0_n77_w133, c0_n77_w134, c0_n77_w135, c0_n77_w136, c0_n77_w137, c0_n77_w138, c0_n77_w139, c0_n77_w140, c0_n77_w141, c0_n77_w142, c0_n77_w143, c0_n77_w144, c0_n77_w145, c0_n77_w146, c0_n77_w147, c0_n77_w148, c0_n77_w149, c0_n77_w150, c0_n77_w151, c0_n77_w152, c0_n77_w153, c0_n77_w154, c0_n77_w155, c0_n77_w156, c0_n77_w157, c0_n77_w158, c0_n77_w159, c0_n77_w160, c0_n77_w161, c0_n77_w162, c0_n77_w163, c0_n77_w164, c0_n77_w165, c0_n77_w166, c0_n77_w167, c0_n77_w168, c0_n77_w169, c0_n77_w170, c0_n77_w171, c0_n77_w172, c0_n77_w173, c0_n77_w174, c0_n77_w175, c0_n77_w176, c0_n77_w177, c0_n77_w178, c0_n77_w179, c0_n77_w180, c0_n77_w181, c0_n77_w182, c0_n77_w183, c0_n77_w184, c0_n77_w185, c0_n77_w186, c0_n77_w187, c0_n77_w188, c0_n77_w189, c0_n77_w190, c0_n77_w191, c0_n77_w192, c0_n77_w193, c0_n77_w194, c0_n77_w195, c0_n77_w196, c0_n77_w197, c0_n77_w198, c0_n77_w199, c0_n77_w200, c0_n78_w1, c0_n78_w2, c0_n78_w3, c0_n78_w4, c0_n78_w5, c0_n78_w6, c0_n78_w7, c0_n78_w8, c0_n78_w9, c0_n78_w10, c0_n78_w11, c0_n78_w12, c0_n78_w13, c0_n78_w14, c0_n78_w15, c0_n78_w16, c0_n78_w17, c0_n78_w18, c0_n78_w19, c0_n78_w20, c0_n78_w21, c0_n78_w22, c0_n78_w23, c0_n78_w24, c0_n78_w25, c0_n78_w26, c0_n78_w27, c0_n78_w28, c0_n78_w29, c0_n78_w30, c0_n78_w31, c0_n78_w32, c0_n78_w33, c0_n78_w34, c0_n78_w35, c0_n78_w36, c0_n78_w37, c0_n78_w38, c0_n78_w39, c0_n78_w40, c0_n78_w41, c0_n78_w42, c0_n78_w43, c0_n78_w44, c0_n78_w45, c0_n78_w46, c0_n78_w47, c0_n78_w48, c0_n78_w49, c0_n78_w50, c0_n78_w51, c0_n78_w52, c0_n78_w53, c0_n78_w54, c0_n78_w55, c0_n78_w56, c0_n78_w57, c0_n78_w58, c0_n78_w59, c0_n78_w60, c0_n78_w61, c0_n78_w62, c0_n78_w63, c0_n78_w64, c0_n78_w65, c0_n78_w66, c0_n78_w67, c0_n78_w68, c0_n78_w69, c0_n78_w70, c0_n78_w71, c0_n78_w72, c0_n78_w73, c0_n78_w74, c0_n78_w75, c0_n78_w76, c0_n78_w77, c0_n78_w78, c0_n78_w79, c0_n78_w80, c0_n78_w81, c0_n78_w82, c0_n78_w83, c0_n78_w84, c0_n78_w85, c0_n78_w86, c0_n78_w87, c0_n78_w88, c0_n78_w89, c0_n78_w90, c0_n78_w91, c0_n78_w92, c0_n78_w93, c0_n78_w94, c0_n78_w95, c0_n78_w96, c0_n78_w97, c0_n78_w98, c0_n78_w99, c0_n78_w100, c0_n78_w101, c0_n78_w102, c0_n78_w103, c0_n78_w104, c0_n78_w105, c0_n78_w106, c0_n78_w107, c0_n78_w108, c0_n78_w109, c0_n78_w110, c0_n78_w111, c0_n78_w112, c0_n78_w113, c0_n78_w114, c0_n78_w115, c0_n78_w116, c0_n78_w117, c0_n78_w118, c0_n78_w119, c0_n78_w120, c0_n78_w121, c0_n78_w122, c0_n78_w123, c0_n78_w124, c0_n78_w125, c0_n78_w126, c0_n78_w127, c0_n78_w128, c0_n78_w129, c0_n78_w130, c0_n78_w131, c0_n78_w132, c0_n78_w133, c0_n78_w134, c0_n78_w135, c0_n78_w136, c0_n78_w137, c0_n78_w138, c0_n78_w139, c0_n78_w140, c0_n78_w141, c0_n78_w142, c0_n78_w143, c0_n78_w144, c0_n78_w145, c0_n78_w146, c0_n78_w147, c0_n78_w148, c0_n78_w149, c0_n78_w150, c0_n78_w151, c0_n78_w152, c0_n78_w153, c0_n78_w154, c0_n78_w155, c0_n78_w156, c0_n78_w157, c0_n78_w158, c0_n78_w159, c0_n78_w160, c0_n78_w161, c0_n78_w162, c0_n78_w163, c0_n78_w164, c0_n78_w165, c0_n78_w166, c0_n78_w167, c0_n78_w168, c0_n78_w169, c0_n78_w170, c0_n78_w171, c0_n78_w172, c0_n78_w173, c0_n78_w174, c0_n78_w175, c0_n78_w176, c0_n78_w177, c0_n78_w178, c0_n78_w179, c0_n78_w180, c0_n78_w181, c0_n78_w182, c0_n78_w183, c0_n78_w184, c0_n78_w185, c0_n78_w186, c0_n78_w187, c0_n78_w188, c0_n78_w189, c0_n78_w190, c0_n78_w191, c0_n78_w192, c0_n78_w193, c0_n78_w194, c0_n78_w195, c0_n78_w196, c0_n78_w197, c0_n78_w198, c0_n78_w199, c0_n78_w200, c0_n79_w1, c0_n79_w2, c0_n79_w3, c0_n79_w4, c0_n79_w5, c0_n79_w6, c0_n79_w7, c0_n79_w8, c0_n79_w9, c0_n79_w10, c0_n79_w11, c0_n79_w12, c0_n79_w13, c0_n79_w14, c0_n79_w15, c0_n79_w16, c0_n79_w17, c0_n79_w18, c0_n79_w19, c0_n79_w20, c0_n79_w21, c0_n79_w22, c0_n79_w23, c0_n79_w24, c0_n79_w25, c0_n79_w26, c0_n79_w27, c0_n79_w28, c0_n79_w29, c0_n79_w30, c0_n79_w31, c0_n79_w32, c0_n79_w33, c0_n79_w34, c0_n79_w35, c0_n79_w36, c0_n79_w37, c0_n79_w38, c0_n79_w39, c0_n79_w40, c0_n79_w41, c0_n79_w42, c0_n79_w43, c0_n79_w44, c0_n79_w45, c0_n79_w46, c0_n79_w47, c0_n79_w48, c0_n79_w49, c0_n79_w50, c0_n79_w51, c0_n79_w52, c0_n79_w53, c0_n79_w54, c0_n79_w55, c0_n79_w56, c0_n79_w57, c0_n79_w58, c0_n79_w59, c0_n79_w60, c0_n79_w61, c0_n79_w62, c0_n79_w63, c0_n79_w64, c0_n79_w65, c0_n79_w66, c0_n79_w67, c0_n79_w68, c0_n79_w69, c0_n79_w70, c0_n79_w71, c0_n79_w72, c0_n79_w73, c0_n79_w74, c0_n79_w75, c0_n79_w76, c0_n79_w77, c0_n79_w78, c0_n79_w79, c0_n79_w80, c0_n79_w81, c0_n79_w82, c0_n79_w83, c0_n79_w84, c0_n79_w85, c0_n79_w86, c0_n79_w87, c0_n79_w88, c0_n79_w89, c0_n79_w90, c0_n79_w91, c0_n79_w92, c0_n79_w93, c0_n79_w94, c0_n79_w95, c0_n79_w96, c0_n79_w97, c0_n79_w98, c0_n79_w99, c0_n79_w100, c0_n79_w101, c0_n79_w102, c0_n79_w103, c0_n79_w104, c0_n79_w105, c0_n79_w106, c0_n79_w107, c0_n79_w108, c0_n79_w109, c0_n79_w110, c0_n79_w111, c0_n79_w112, c0_n79_w113, c0_n79_w114, c0_n79_w115, c0_n79_w116, c0_n79_w117, c0_n79_w118, c0_n79_w119, c0_n79_w120, c0_n79_w121, c0_n79_w122, c0_n79_w123, c0_n79_w124, c0_n79_w125, c0_n79_w126, c0_n79_w127, c0_n79_w128, c0_n79_w129, c0_n79_w130, c0_n79_w131, c0_n79_w132, c0_n79_w133, c0_n79_w134, c0_n79_w135, c0_n79_w136, c0_n79_w137, c0_n79_w138, c0_n79_w139, c0_n79_w140, c0_n79_w141, c0_n79_w142, c0_n79_w143, c0_n79_w144, c0_n79_w145, c0_n79_w146, c0_n79_w147, c0_n79_w148, c0_n79_w149, c0_n79_w150, c0_n79_w151, c0_n79_w152, c0_n79_w153, c0_n79_w154, c0_n79_w155, c0_n79_w156, c0_n79_w157, c0_n79_w158, c0_n79_w159, c0_n79_w160, c0_n79_w161, c0_n79_w162, c0_n79_w163, c0_n79_w164, c0_n79_w165, c0_n79_w166, c0_n79_w167, c0_n79_w168, c0_n79_w169, c0_n79_w170, c0_n79_w171, c0_n79_w172, c0_n79_w173, c0_n79_w174, c0_n79_w175, c0_n79_w176, c0_n79_w177, c0_n79_w178, c0_n79_w179, c0_n79_w180, c0_n79_w181, c0_n79_w182, c0_n79_w183, c0_n79_w184, c0_n79_w185, c0_n79_w186, c0_n79_w187, c0_n79_w188, c0_n79_w189, c0_n79_w190, c0_n79_w191, c0_n79_w192, c0_n79_w193, c0_n79_w194, c0_n79_w195, c0_n79_w196, c0_n79_w197, c0_n79_w198, c0_n79_w199, c0_n79_w200, c0_n80_w1, c0_n80_w2, c0_n80_w3, c0_n80_w4, c0_n80_w5, c0_n80_w6, c0_n80_w7, c0_n80_w8, c0_n80_w9, c0_n80_w10, c0_n80_w11, c0_n80_w12, c0_n80_w13, c0_n80_w14, c0_n80_w15, c0_n80_w16, c0_n80_w17, c0_n80_w18, c0_n80_w19, c0_n80_w20, c0_n80_w21, c0_n80_w22, c0_n80_w23, c0_n80_w24, c0_n80_w25, c0_n80_w26, c0_n80_w27, c0_n80_w28, c0_n80_w29, c0_n80_w30, c0_n80_w31, c0_n80_w32, c0_n80_w33, c0_n80_w34, c0_n80_w35, c0_n80_w36, c0_n80_w37, c0_n80_w38, c0_n80_w39, c0_n80_w40, c0_n80_w41, c0_n80_w42, c0_n80_w43, c0_n80_w44, c0_n80_w45, c0_n80_w46, c0_n80_w47, c0_n80_w48, c0_n80_w49, c0_n80_w50, c0_n80_w51, c0_n80_w52, c0_n80_w53, c0_n80_w54, c0_n80_w55, c0_n80_w56, c0_n80_w57, c0_n80_w58, c0_n80_w59, c0_n80_w60, c0_n80_w61, c0_n80_w62, c0_n80_w63, c0_n80_w64, c0_n80_w65, c0_n80_w66, c0_n80_w67, c0_n80_w68, c0_n80_w69, c0_n80_w70, c0_n80_w71, c0_n80_w72, c0_n80_w73, c0_n80_w74, c0_n80_w75, c0_n80_w76, c0_n80_w77, c0_n80_w78, c0_n80_w79, c0_n80_w80, c0_n80_w81, c0_n80_w82, c0_n80_w83, c0_n80_w84, c0_n80_w85, c0_n80_w86, c0_n80_w87, c0_n80_w88, c0_n80_w89, c0_n80_w90, c0_n80_w91, c0_n80_w92, c0_n80_w93, c0_n80_w94, c0_n80_w95, c0_n80_w96, c0_n80_w97, c0_n80_w98, c0_n80_w99, c0_n80_w100, c0_n80_w101, c0_n80_w102, c0_n80_w103, c0_n80_w104, c0_n80_w105, c0_n80_w106, c0_n80_w107, c0_n80_w108, c0_n80_w109, c0_n80_w110, c0_n80_w111, c0_n80_w112, c0_n80_w113, c0_n80_w114, c0_n80_w115, c0_n80_w116, c0_n80_w117, c0_n80_w118, c0_n80_w119, c0_n80_w120, c0_n80_w121, c0_n80_w122, c0_n80_w123, c0_n80_w124, c0_n80_w125, c0_n80_w126, c0_n80_w127, c0_n80_w128, c0_n80_w129, c0_n80_w130, c0_n80_w131, c0_n80_w132, c0_n80_w133, c0_n80_w134, c0_n80_w135, c0_n80_w136, c0_n80_w137, c0_n80_w138, c0_n80_w139, c0_n80_w140, c0_n80_w141, c0_n80_w142, c0_n80_w143, c0_n80_w144, c0_n80_w145, c0_n80_w146, c0_n80_w147, c0_n80_w148, c0_n80_w149, c0_n80_w150, c0_n80_w151, c0_n80_w152, c0_n80_w153, c0_n80_w154, c0_n80_w155, c0_n80_w156, c0_n80_w157, c0_n80_w158, c0_n80_w159, c0_n80_w160, c0_n80_w161, c0_n80_w162, c0_n80_w163, c0_n80_w164, c0_n80_w165, c0_n80_w166, c0_n80_w167, c0_n80_w168, c0_n80_w169, c0_n80_w170, c0_n80_w171, c0_n80_w172, c0_n80_w173, c0_n80_w174, c0_n80_w175, c0_n80_w176, c0_n80_w177, c0_n80_w178, c0_n80_w179, c0_n80_w180, c0_n80_w181, c0_n80_w182, c0_n80_w183, c0_n80_w184, c0_n80_w185, c0_n80_w186, c0_n80_w187, c0_n80_w188, c0_n80_w189, c0_n80_w190, c0_n80_w191, c0_n80_w192, c0_n80_w193, c0_n80_w194, c0_n80_w195, c0_n80_w196, c0_n80_w197, c0_n80_w198, c0_n80_w199, c0_n80_w200, c0_n81_w1, c0_n81_w2, c0_n81_w3, c0_n81_w4, c0_n81_w5, c0_n81_w6, c0_n81_w7, c0_n81_w8, c0_n81_w9, c0_n81_w10, c0_n81_w11, c0_n81_w12, c0_n81_w13, c0_n81_w14, c0_n81_w15, c0_n81_w16, c0_n81_w17, c0_n81_w18, c0_n81_w19, c0_n81_w20, c0_n81_w21, c0_n81_w22, c0_n81_w23, c0_n81_w24, c0_n81_w25, c0_n81_w26, c0_n81_w27, c0_n81_w28, c0_n81_w29, c0_n81_w30, c0_n81_w31, c0_n81_w32, c0_n81_w33, c0_n81_w34, c0_n81_w35, c0_n81_w36, c0_n81_w37, c0_n81_w38, c0_n81_w39, c0_n81_w40, c0_n81_w41, c0_n81_w42, c0_n81_w43, c0_n81_w44, c0_n81_w45, c0_n81_w46, c0_n81_w47, c0_n81_w48, c0_n81_w49, c0_n81_w50, c0_n81_w51, c0_n81_w52, c0_n81_w53, c0_n81_w54, c0_n81_w55, c0_n81_w56, c0_n81_w57, c0_n81_w58, c0_n81_w59, c0_n81_w60, c0_n81_w61, c0_n81_w62, c0_n81_w63, c0_n81_w64, c0_n81_w65, c0_n81_w66, c0_n81_w67, c0_n81_w68, c0_n81_w69, c0_n81_w70, c0_n81_w71, c0_n81_w72, c0_n81_w73, c0_n81_w74, c0_n81_w75, c0_n81_w76, c0_n81_w77, c0_n81_w78, c0_n81_w79, c0_n81_w80, c0_n81_w81, c0_n81_w82, c0_n81_w83, c0_n81_w84, c0_n81_w85, c0_n81_w86, c0_n81_w87, c0_n81_w88, c0_n81_w89, c0_n81_w90, c0_n81_w91, c0_n81_w92, c0_n81_w93, c0_n81_w94, c0_n81_w95, c0_n81_w96, c0_n81_w97, c0_n81_w98, c0_n81_w99, c0_n81_w100, c0_n81_w101, c0_n81_w102, c0_n81_w103, c0_n81_w104, c0_n81_w105, c0_n81_w106, c0_n81_w107, c0_n81_w108, c0_n81_w109, c0_n81_w110, c0_n81_w111, c0_n81_w112, c0_n81_w113, c0_n81_w114, c0_n81_w115, c0_n81_w116, c0_n81_w117, c0_n81_w118, c0_n81_w119, c0_n81_w120, c0_n81_w121, c0_n81_w122, c0_n81_w123, c0_n81_w124, c0_n81_w125, c0_n81_w126, c0_n81_w127, c0_n81_w128, c0_n81_w129, c0_n81_w130, c0_n81_w131, c0_n81_w132, c0_n81_w133, c0_n81_w134, c0_n81_w135, c0_n81_w136, c0_n81_w137, c0_n81_w138, c0_n81_w139, c0_n81_w140, c0_n81_w141, c0_n81_w142, c0_n81_w143, c0_n81_w144, c0_n81_w145, c0_n81_w146, c0_n81_w147, c0_n81_w148, c0_n81_w149, c0_n81_w150, c0_n81_w151, c0_n81_w152, c0_n81_w153, c0_n81_w154, c0_n81_w155, c0_n81_w156, c0_n81_w157, c0_n81_w158, c0_n81_w159, c0_n81_w160, c0_n81_w161, c0_n81_w162, c0_n81_w163, c0_n81_w164, c0_n81_w165, c0_n81_w166, c0_n81_w167, c0_n81_w168, c0_n81_w169, c0_n81_w170, c0_n81_w171, c0_n81_w172, c0_n81_w173, c0_n81_w174, c0_n81_w175, c0_n81_w176, c0_n81_w177, c0_n81_w178, c0_n81_w179, c0_n81_w180, c0_n81_w181, c0_n81_w182, c0_n81_w183, c0_n81_w184, c0_n81_w185, c0_n81_w186, c0_n81_w187, c0_n81_w188, c0_n81_w189, c0_n81_w190, c0_n81_w191, c0_n81_w192, c0_n81_w193, c0_n81_w194, c0_n81_w195, c0_n81_w196, c0_n81_w197, c0_n81_w198, c0_n81_w199, c0_n81_w200, c0_n82_w1, c0_n82_w2, c0_n82_w3, c0_n82_w4, c0_n82_w5, c0_n82_w6, c0_n82_w7, c0_n82_w8, c0_n82_w9, c0_n82_w10, c0_n82_w11, c0_n82_w12, c0_n82_w13, c0_n82_w14, c0_n82_w15, c0_n82_w16, c0_n82_w17, c0_n82_w18, c0_n82_w19, c0_n82_w20, c0_n82_w21, c0_n82_w22, c0_n82_w23, c0_n82_w24, c0_n82_w25, c0_n82_w26, c0_n82_w27, c0_n82_w28, c0_n82_w29, c0_n82_w30, c0_n82_w31, c0_n82_w32, c0_n82_w33, c0_n82_w34, c0_n82_w35, c0_n82_w36, c0_n82_w37, c0_n82_w38, c0_n82_w39, c0_n82_w40, c0_n82_w41, c0_n82_w42, c0_n82_w43, c0_n82_w44, c0_n82_w45, c0_n82_w46, c0_n82_w47, c0_n82_w48, c0_n82_w49, c0_n82_w50, c0_n82_w51, c0_n82_w52, c0_n82_w53, c0_n82_w54, c0_n82_w55, c0_n82_w56, c0_n82_w57, c0_n82_w58, c0_n82_w59, c0_n82_w60, c0_n82_w61, c0_n82_w62, c0_n82_w63, c0_n82_w64, c0_n82_w65, c0_n82_w66, c0_n82_w67, c0_n82_w68, c0_n82_w69, c0_n82_w70, c0_n82_w71, c0_n82_w72, c0_n82_w73, c0_n82_w74, c0_n82_w75, c0_n82_w76, c0_n82_w77, c0_n82_w78, c0_n82_w79, c0_n82_w80, c0_n82_w81, c0_n82_w82, c0_n82_w83, c0_n82_w84, c0_n82_w85, c0_n82_w86, c0_n82_w87, c0_n82_w88, c0_n82_w89, c0_n82_w90, c0_n82_w91, c0_n82_w92, c0_n82_w93, c0_n82_w94, c0_n82_w95, c0_n82_w96, c0_n82_w97, c0_n82_w98, c0_n82_w99, c0_n82_w100, c0_n82_w101, c0_n82_w102, c0_n82_w103, c0_n82_w104, c0_n82_w105, c0_n82_w106, c0_n82_w107, c0_n82_w108, c0_n82_w109, c0_n82_w110, c0_n82_w111, c0_n82_w112, c0_n82_w113, c0_n82_w114, c0_n82_w115, c0_n82_w116, c0_n82_w117, c0_n82_w118, c0_n82_w119, c0_n82_w120, c0_n82_w121, c0_n82_w122, c0_n82_w123, c0_n82_w124, c0_n82_w125, c0_n82_w126, c0_n82_w127, c0_n82_w128, c0_n82_w129, c0_n82_w130, c0_n82_w131, c0_n82_w132, c0_n82_w133, c0_n82_w134, c0_n82_w135, c0_n82_w136, c0_n82_w137, c0_n82_w138, c0_n82_w139, c0_n82_w140, c0_n82_w141, c0_n82_w142, c0_n82_w143, c0_n82_w144, c0_n82_w145, c0_n82_w146, c0_n82_w147, c0_n82_w148, c0_n82_w149, c0_n82_w150, c0_n82_w151, c0_n82_w152, c0_n82_w153, c0_n82_w154, c0_n82_w155, c0_n82_w156, c0_n82_w157, c0_n82_w158, c0_n82_w159, c0_n82_w160, c0_n82_w161, c0_n82_w162, c0_n82_w163, c0_n82_w164, c0_n82_w165, c0_n82_w166, c0_n82_w167, c0_n82_w168, c0_n82_w169, c0_n82_w170, c0_n82_w171, c0_n82_w172, c0_n82_w173, c0_n82_w174, c0_n82_w175, c0_n82_w176, c0_n82_w177, c0_n82_w178, c0_n82_w179, c0_n82_w180, c0_n82_w181, c0_n82_w182, c0_n82_w183, c0_n82_w184, c0_n82_w185, c0_n82_w186, c0_n82_w187, c0_n82_w188, c0_n82_w189, c0_n82_w190, c0_n82_w191, c0_n82_w192, c0_n82_w193, c0_n82_w194, c0_n82_w195, c0_n82_w196, c0_n82_w197, c0_n82_w198, c0_n82_w199, c0_n82_w200, c0_n83_w1, c0_n83_w2, c0_n83_w3, c0_n83_w4, c0_n83_w5, c0_n83_w6, c0_n83_w7, c0_n83_w8, c0_n83_w9, c0_n83_w10, c0_n83_w11, c0_n83_w12, c0_n83_w13, c0_n83_w14, c0_n83_w15, c0_n83_w16, c0_n83_w17, c0_n83_w18, c0_n83_w19, c0_n83_w20, c0_n83_w21, c0_n83_w22, c0_n83_w23, c0_n83_w24, c0_n83_w25, c0_n83_w26, c0_n83_w27, c0_n83_w28, c0_n83_w29, c0_n83_w30, c0_n83_w31, c0_n83_w32, c0_n83_w33, c0_n83_w34, c0_n83_w35, c0_n83_w36, c0_n83_w37, c0_n83_w38, c0_n83_w39, c0_n83_w40, c0_n83_w41, c0_n83_w42, c0_n83_w43, c0_n83_w44, c0_n83_w45, c0_n83_w46, c0_n83_w47, c0_n83_w48, c0_n83_w49, c0_n83_w50, c0_n83_w51, c0_n83_w52, c0_n83_w53, c0_n83_w54, c0_n83_w55, c0_n83_w56, c0_n83_w57, c0_n83_w58, c0_n83_w59, c0_n83_w60, c0_n83_w61, c0_n83_w62, c0_n83_w63, c0_n83_w64, c0_n83_w65, c0_n83_w66, c0_n83_w67, c0_n83_w68, c0_n83_w69, c0_n83_w70, c0_n83_w71, c0_n83_w72, c0_n83_w73, c0_n83_w74, c0_n83_w75, c0_n83_w76, c0_n83_w77, c0_n83_w78, c0_n83_w79, c0_n83_w80, c0_n83_w81, c0_n83_w82, c0_n83_w83, c0_n83_w84, c0_n83_w85, c0_n83_w86, c0_n83_w87, c0_n83_w88, c0_n83_w89, c0_n83_w90, c0_n83_w91, c0_n83_w92, c0_n83_w93, c0_n83_w94, c0_n83_w95, c0_n83_w96, c0_n83_w97, c0_n83_w98, c0_n83_w99, c0_n83_w100, c0_n83_w101, c0_n83_w102, c0_n83_w103, c0_n83_w104, c0_n83_w105, c0_n83_w106, c0_n83_w107, c0_n83_w108, c0_n83_w109, c0_n83_w110, c0_n83_w111, c0_n83_w112, c0_n83_w113, c0_n83_w114, c0_n83_w115, c0_n83_w116, c0_n83_w117, c0_n83_w118, c0_n83_w119, c0_n83_w120, c0_n83_w121, c0_n83_w122, c0_n83_w123, c0_n83_w124, c0_n83_w125, c0_n83_w126, c0_n83_w127, c0_n83_w128, c0_n83_w129, c0_n83_w130, c0_n83_w131, c0_n83_w132, c0_n83_w133, c0_n83_w134, c0_n83_w135, c0_n83_w136, c0_n83_w137, c0_n83_w138, c0_n83_w139, c0_n83_w140, c0_n83_w141, c0_n83_w142, c0_n83_w143, c0_n83_w144, c0_n83_w145, c0_n83_w146, c0_n83_w147, c0_n83_w148, c0_n83_w149, c0_n83_w150, c0_n83_w151, c0_n83_w152, c0_n83_w153, c0_n83_w154, c0_n83_w155, c0_n83_w156, c0_n83_w157, c0_n83_w158, c0_n83_w159, c0_n83_w160, c0_n83_w161, c0_n83_w162, c0_n83_w163, c0_n83_w164, c0_n83_w165, c0_n83_w166, c0_n83_w167, c0_n83_w168, c0_n83_w169, c0_n83_w170, c0_n83_w171, c0_n83_w172, c0_n83_w173, c0_n83_w174, c0_n83_w175, c0_n83_w176, c0_n83_w177, c0_n83_w178, c0_n83_w179, c0_n83_w180, c0_n83_w181, c0_n83_w182, c0_n83_w183, c0_n83_w184, c0_n83_w185, c0_n83_w186, c0_n83_w187, c0_n83_w188, c0_n83_w189, c0_n83_w190, c0_n83_w191, c0_n83_w192, c0_n83_w193, c0_n83_w194, c0_n83_w195, c0_n83_w196, c0_n83_w197, c0_n83_w198, c0_n83_w199, c0_n83_w200, c0_n84_w1, c0_n84_w2, c0_n84_w3, c0_n84_w4, c0_n84_w5, c0_n84_w6, c0_n84_w7, c0_n84_w8, c0_n84_w9, c0_n84_w10, c0_n84_w11, c0_n84_w12, c0_n84_w13, c0_n84_w14, c0_n84_w15, c0_n84_w16, c0_n84_w17, c0_n84_w18, c0_n84_w19, c0_n84_w20, c0_n84_w21, c0_n84_w22, c0_n84_w23, c0_n84_w24, c0_n84_w25, c0_n84_w26, c0_n84_w27, c0_n84_w28, c0_n84_w29, c0_n84_w30, c0_n84_w31, c0_n84_w32, c0_n84_w33, c0_n84_w34, c0_n84_w35, c0_n84_w36, c0_n84_w37, c0_n84_w38, c0_n84_w39, c0_n84_w40, c0_n84_w41, c0_n84_w42, c0_n84_w43, c0_n84_w44, c0_n84_w45, c0_n84_w46, c0_n84_w47, c0_n84_w48, c0_n84_w49, c0_n84_w50, c0_n84_w51, c0_n84_w52, c0_n84_w53, c0_n84_w54, c0_n84_w55, c0_n84_w56, c0_n84_w57, c0_n84_w58, c0_n84_w59, c0_n84_w60, c0_n84_w61, c0_n84_w62, c0_n84_w63, c0_n84_w64, c0_n84_w65, c0_n84_w66, c0_n84_w67, c0_n84_w68, c0_n84_w69, c0_n84_w70, c0_n84_w71, c0_n84_w72, c0_n84_w73, c0_n84_w74, c0_n84_w75, c0_n84_w76, c0_n84_w77, c0_n84_w78, c0_n84_w79, c0_n84_w80, c0_n84_w81, c0_n84_w82, c0_n84_w83, c0_n84_w84, c0_n84_w85, c0_n84_w86, c0_n84_w87, c0_n84_w88, c0_n84_w89, c0_n84_w90, c0_n84_w91, c0_n84_w92, c0_n84_w93, c0_n84_w94, c0_n84_w95, c0_n84_w96, c0_n84_w97, c0_n84_w98, c0_n84_w99, c0_n84_w100, c0_n84_w101, c0_n84_w102, c0_n84_w103, c0_n84_w104, c0_n84_w105, c0_n84_w106, c0_n84_w107, c0_n84_w108, c0_n84_w109, c0_n84_w110, c0_n84_w111, c0_n84_w112, c0_n84_w113, c0_n84_w114, c0_n84_w115, c0_n84_w116, c0_n84_w117, c0_n84_w118, c0_n84_w119, c0_n84_w120, c0_n84_w121, c0_n84_w122, c0_n84_w123, c0_n84_w124, c0_n84_w125, c0_n84_w126, c0_n84_w127, c0_n84_w128, c0_n84_w129, c0_n84_w130, c0_n84_w131, c0_n84_w132, c0_n84_w133, c0_n84_w134, c0_n84_w135, c0_n84_w136, c0_n84_w137, c0_n84_w138, c0_n84_w139, c0_n84_w140, c0_n84_w141, c0_n84_w142, c0_n84_w143, c0_n84_w144, c0_n84_w145, c0_n84_w146, c0_n84_w147, c0_n84_w148, c0_n84_w149, c0_n84_w150, c0_n84_w151, c0_n84_w152, c0_n84_w153, c0_n84_w154, c0_n84_w155, c0_n84_w156, c0_n84_w157, c0_n84_w158, c0_n84_w159, c0_n84_w160, c0_n84_w161, c0_n84_w162, c0_n84_w163, c0_n84_w164, c0_n84_w165, c0_n84_w166, c0_n84_w167, c0_n84_w168, c0_n84_w169, c0_n84_w170, c0_n84_w171, c0_n84_w172, c0_n84_w173, c0_n84_w174, c0_n84_w175, c0_n84_w176, c0_n84_w177, c0_n84_w178, c0_n84_w179, c0_n84_w180, c0_n84_w181, c0_n84_w182, c0_n84_w183, c0_n84_w184, c0_n84_w185, c0_n84_w186, c0_n84_w187, c0_n84_w188, c0_n84_w189, c0_n84_w190, c0_n84_w191, c0_n84_w192, c0_n84_w193, c0_n84_w194, c0_n84_w195, c0_n84_w196, c0_n84_w197, c0_n84_w198, c0_n84_w199, c0_n84_w200, c0_n85_w1, c0_n85_w2, c0_n85_w3, c0_n85_w4, c0_n85_w5, c0_n85_w6, c0_n85_w7, c0_n85_w8, c0_n85_w9, c0_n85_w10, c0_n85_w11, c0_n85_w12, c0_n85_w13, c0_n85_w14, c0_n85_w15, c0_n85_w16, c0_n85_w17, c0_n85_w18, c0_n85_w19, c0_n85_w20, c0_n85_w21, c0_n85_w22, c0_n85_w23, c0_n85_w24, c0_n85_w25, c0_n85_w26, c0_n85_w27, c0_n85_w28, c0_n85_w29, c0_n85_w30, c0_n85_w31, c0_n85_w32, c0_n85_w33, c0_n85_w34, c0_n85_w35, c0_n85_w36, c0_n85_w37, c0_n85_w38, c0_n85_w39, c0_n85_w40, c0_n85_w41, c0_n85_w42, c0_n85_w43, c0_n85_w44, c0_n85_w45, c0_n85_w46, c0_n85_w47, c0_n85_w48, c0_n85_w49, c0_n85_w50, c0_n85_w51, c0_n85_w52, c0_n85_w53, c0_n85_w54, c0_n85_w55, c0_n85_w56, c0_n85_w57, c0_n85_w58, c0_n85_w59, c0_n85_w60, c0_n85_w61, c0_n85_w62, c0_n85_w63, c0_n85_w64, c0_n85_w65, c0_n85_w66, c0_n85_w67, c0_n85_w68, c0_n85_w69, c0_n85_w70, c0_n85_w71, c0_n85_w72, c0_n85_w73, c0_n85_w74, c0_n85_w75, c0_n85_w76, c0_n85_w77, c0_n85_w78, c0_n85_w79, c0_n85_w80, c0_n85_w81, c0_n85_w82, c0_n85_w83, c0_n85_w84, c0_n85_w85, c0_n85_w86, c0_n85_w87, c0_n85_w88, c0_n85_w89, c0_n85_w90, c0_n85_w91, c0_n85_w92, c0_n85_w93, c0_n85_w94, c0_n85_w95, c0_n85_w96, c0_n85_w97, c0_n85_w98, c0_n85_w99, c0_n85_w100, c0_n85_w101, c0_n85_w102, c0_n85_w103, c0_n85_w104, c0_n85_w105, c0_n85_w106, c0_n85_w107, c0_n85_w108, c0_n85_w109, c0_n85_w110, c0_n85_w111, c0_n85_w112, c0_n85_w113, c0_n85_w114, c0_n85_w115, c0_n85_w116, c0_n85_w117, c0_n85_w118, c0_n85_w119, c0_n85_w120, c0_n85_w121, c0_n85_w122, c0_n85_w123, c0_n85_w124, c0_n85_w125, c0_n85_w126, c0_n85_w127, c0_n85_w128, c0_n85_w129, c0_n85_w130, c0_n85_w131, c0_n85_w132, c0_n85_w133, c0_n85_w134, c0_n85_w135, c0_n85_w136, c0_n85_w137, c0_n85_w138, c0_n85_w139, c0_n85_w140, c0_n85_w141, c0_n85_w142, c0_n85_w143, c0_n85_w144, c0_n85_w145, c0_n85_w146, c0_n85_w147, c0_n85_w148, c0_n85_w149, c0_n85_w150, c0_n85_w151, c0_n85_w152, c0_n85_w153, c0_n85_w154, c0_n85_w155, c0_n85_w156, c0_n85_w157, c0_n85_w158, c0_n85_w159, c0_n85_w160, c0_n85_w161, c0_n85_w162, c0_n85_w163, c0_n85_w164, c0_n85_w165, c0_n85_w166, c0_n85_w167, c0_n85_w168, c0_n85_w169, c0_n85_w170, c0_n85_w171, c0_n85_w172, c0_n85_w173, c0_n85_w174, c0_n85_w175, c0_n85_w176, c0_n85_w177, c0_n85_w178, c0_n85_w179, c0_n85_w180, c0_n85_w181, c0_n85_w182, c0_n85_w183, c0_n85_w184, c0_n85_w185, c0_n85_w186, c0_n85_w187, c0_n85_w188, c0_n85_w189, c0_n85_w190, c0_n85_w191, c0_n85_w192, c0_n85_w193, c0_n85_w194, c0_n85_w195, c0_n85_w196, c0_n85_w197, c0_n85_w198, c0_n85_w199, c0_n85_w200, c0_n86_w1, c0_n86_w2, c0_n86_w3, c0_n86_w4, c0_n86_w5, c0_n86_w6, c0_n86_w7, c0_n86_w8, c0_n86_w9, c0_n86_w10, c0_n86_w11, c0_n86_w12, c0_n86_w13, c0_n86_w14, c0_n86_w15, c0_n86_w16, c0_n86_w17, c0_n86_w18, c0_n86_w19, c0_n86_w20, c0_n86_w21, c0_n86_w22, c0_n86_w23, c0_n86_w24, c0_n86_w25, c0_n86_w26, c0_n86_w27, c0_n86_w28, c0_n86_w29, c0_n86_w30, c0_n86_w31, c0_n86_w32, c0_n86_w33, c0_n86_w34, c0_n86_w35, c0_n86_w36, c0_n86_w37, c0_n86_w38, c0_n86_w39, c0_n86_w40, c0_n86_w41, c0_n86_w42, c0_n86_w43, c0_n86_w44, c0_n86_w45, c0_n86_w46, c0_n86_w47, c0_n86_w48, c0_n86_w49, c0_n86_w50, c0_n86_w51, c0_n86_w52, c0_n86_w53, c0_n86_w54, c0_n86_w55, c0_n86_w56, c0_n86_w57, c0_n86_w58, c0_n86_w59, c0_n86_w60, c0_n86_w61, c0_n86_w62, c0_n86_w63, c0_n86_w64, c0_n86_w65, c0_n86_w66, c0_n86_w67, c0_n86_w68, c0_n86_w69, c0_n86_w70, c0_n86_w71, c0_n86_w72, c0_n86_w73, c0_n86_w74, c0_n86_w75, c0_n86_w76, c0_n86_w77, c0_n86_w78, c0_n86_w79, c0_n86_w80, c0_n86_w81, c0_n86_w82, c0_n86_w83, c0_n86_w84, c0_n86_w85, c0_n86_w86, c0_n86_w87, c0_n86_w88, c0_n86_w89, c0_n86_w90, c0_n86_w91, c0_n86_w92, c0_n86_w93, c0_n86_w94, c0_n86_w95, c0_n86_w96, c0_n86_w97, c0_n86_w98, c0_n86_w99, c0_n86_w100, c0_n86_w101, c0_n86_w102, c0_n86_w103, c0_n86_w104, c0_n86_w105, c0_n86_w106, c0_n86_w107, c0_n86_w108, c0_n86_w109, c0_n86_w110, c0_n86_w111, c0_n86_w112, c0_n86_w113, c0_n86_w114, c0_n86_w115, c0_n86_w116, c0_n86_w117, c0_n86_w118, c0_n86_w119, c0_n86_w120, c0_n86_w121, c0_n86_w122, c0_n86_w123, c0_n86_w124, c0_n86_w125, c0_n86_w126, c0_n86_w127, c0_n86_w128, c0_n86_w129, c0_n86_w130, c0_n86_w131, c0_n86_w132, c0_n86_w133, c0_n86_w134, c0_n86_w135, c0_n86_w136, c0_n86_w137, c0_n86_w138, c0_n86_w139, c0_n86_w140, c0_n86_w141, c0_n86_w142, c0_n86_w143, c0_n86_w144, c0_n86_w145, c0_n86_w146, c0_n86_w147, c0_n86_w148, c0_n86_w149, c0_n86_w150, c0_n86_w151, c0_n86_w152, c0_n86_w153, c0_n86_w154, c0_n86_w155, c0_n86_w156, c0_n86_w157, c0_n86_w158, c0_n86_w159, c0_n86_w160, c0_n86_w161, c0_n86_w162, c0_n86_w163, c0_n86_w164, c0_n86_w165, c0_n86_w166, c0_n86_w167, c0_n86_w168, c0_n86_w169, c0_n86_w170, c0_n86_w171, c0_n86_w172, c0_n86_w173, c0_n86_w174, c0_n86_w175, c0_n86_w176, c0_n86_w177, c0_n86_w178, c0_n86_w179, c0_n86_w180, c0_n86_w181, c0_n86_w182, c0_n86_w183, c0_n86_w184, c0_n86_w185, c0_n86_w186, c0_n86_w187, c0_n86_w188, c0_n86_w189, c0_n86_w190, c0_n86_w191, c0_n86_w192, c0_n86_w193, c0_n86_w194, c0_n86_w195, c0_n86_w196, c0_n86_w197, c0_n86_w198, c0_n86_w199, c0_n86_w200, c0_n87_w1, c0_n87_w2, c0_n87_w3, c0_n87_w4, c0_n87_w5, c0_n87_w6, c0_n87_w7, c0_n87_w8, c0_n87_w9, c0_n87_w10, c0_n87_w11, c0_n87_w12, c0_n87_w13, c0_n87_w14, c0_n87_w15, c0_n87_w16, c0_n87_w17, c0_n87_w18, c0_n87_w19, c0_n87_w20, c0_n87_w21, c0_n87_w22, c0_n87_w23, c0_n87_w24, c0_n87_w25, c0_n87_w26, c0_n87_w27, c0_n87_w28, c0_n87_w29, c0_n87_w30, c0_n87_w31, c0_n87_w32, c0_n87_w33, c0_n87_w34, c0_n87_w35, c0_n87_w36, c0_n87_w37, c0_n87_w38, c0_n87_w39, c0_n87_w40, c0_n87_w41, c0_n87_w42, c0_n87_w43, c0_n87_w44, c0_n87_w45, c0_n87_w46, c0_n87_w47, c0_n87_w48, c0_n87_w49, c0_n87_w50, c0_n87_w51, c0_n87_w52, c0_n87_w53, c0_n87_w54, c0_n87_w55, c0_n87_w56, c0_n87_w57, c0_n87_w58, c0_n87_w59, c0_n87_w60, c0_n87_w61, c0_n87_w62, c0_n87_w63, c0_n87_w64, c0_n87_w65, c0_n87_w66, c0_n87_w67, c0_n87_w68, c0_n87_w69, c0_n87_w70, c0_n87_w71, c0_n87_w72, c0_n87_w73, c0_n87_w74, c0_n87_w75, c0_n87_w76, c0_n87_w77, c0_n87_w78, c0_n87_w79, c0_n87_w80, c0_n87_w81, c0_n87_w82, c0_n87_w83, c0_n87_w84, c0_n87_w85, c0_n87_w86, c0_n87_w87, c0_n87_w88, c0_n87_w89, c0_n87_w90, c0_n87_w91, c0_n87_w92, c0_n87_w93, c0_n87_w94, c0_n87_w95, c0_n87_w96, c0_n87_w97, c0_n87_w98, c0_n87_w99, c0_n87_w100, c0_n87_w101, c0_n87_w102, c0_n87_w103, c0_n87_w104, c0_n87_w105, c0_n87_w106, c0_n87_w107, c0_n87_w108, c0_n87_w109, c0_n87_w110, c0_n87_w111, c0_n87_w112, c0_n87_w113, c0_n87_w114, c0_n87_w115, c0_n87_w116, c0_n87_w117, c0_n87_w118, c0_n87_w119, c0_n87_w120, c0_n87_w121, c0_n87_w122, c0_n87_w123, c0_n87_w124, c0_n87_w125, c0_n87_w126, c0_n87_w127, c0_n87_w128, c0_n87_w129, c0_n87_w130, c0_n87_w131, c0_n87_w132, c0_n87_w133, c0_n87_w134, c0_n87_w135, c0_n87_w136, c0_n87_w137, c0_n87_w138, c0_n87_w139, c0_n87_w140, c0_n87_w141, c0_n87_w142, c0_n87_w143, c0_n87_w144, c0_n87_w145, c0_n87_w146, c0_n87_w147, c0_n87_w148, c0_n87_w149, c0_n87_w150, c0_n87_w151, c0_n87_w152, c0_n87_w153, c0_n87_w154, c0_n87_w155, c0_n87_w156, c0_n87_w157, c0_n87_w158, c0_n87_w159, c0_n87_w160, c0_n87_w161, c0_n87_w162, c0_n87_w163, c0_n87_w164, c0_n87_w165, c0_n87_w166, c0_n87_w167, c0_n87_w168, c0_n87_w169, c0_n87_w170, c0_n87_w171, c0_n87_w172, c0_n87_w173, c0_n87_w174, c0_n87_w175, c0_n87_w176, c0_n87_w177, c0_n87_w178, c0_n87_w179, c0_n87_w180, c0_n87_w181, c0_n87_w182, c0_n87_w183, c0_n87_w184, c0_n87_w185, c0_n87_w186, c0_n87_w187, c0_n87_w188, c0_n87_w189, c0_n87_w190, c0_n87_w191, c0_n87_w192, c0_n87_w193, c0_n87_w194, c0_n87_w195, c0_n87_w196, c0_n87_w197, c0_n87_w198, c0_n87_w199, c0_n87_w200, c0_n88_w1, c0_n88_w2, c0_n88_w3, c0_n88_w4, c0_n88_w5, c0_n88_w6, c0_n88_w7, c0_n88_w8, c0_n88_w9, c0_n88_w10, c0_n88_w11, c0_n88_w12, c0_n88_w13, c0_n88_w14, c0_n88_w15, c0_n88_w16, c0_n88_w17, c0_n88_w18, c0_n88_w19, c0_n88_w20, c0_n88_w21, c0_n88_w22, c0_n88_w23, c0_n88_w24, c0_n88_w25, c0_n88_w26, c0_n88_w27, c0_n88_w28, c0_n88_w29, c0_n88_w30, c0_n88_w31, c0_n88_w32, c0_n88_w33, c0_n88_w34, c0_n88_w35, c0_n88_w36, c0_n88_w37, c0_n88_w38, c0_n88_w39, c0_n88_w40, c0_n88_w41, c0_n88_w42, c0_n88_w43, c0_n88_w44, c0_n88_w45, c0_n88_w46, c0_n88_w47, c0_n88_w48, c0_n88_w49, c0_n88_w50, c0_n88_w51, c0_n88_w52, c0_n88_w53, c0_n88_w54, c0_n88_w55, c0_n88_w56, c0_n88_w57, c0_n88_w58, c0_n88_w59, c0_n88_w60, c0_n88_w61, c0_n88_w62, c0_n88_w63, c0_n88_w64, c0_n88_w65, c0_n88_w66, c0_n88_w67, c0_n88_w68, c0_n88_w69, c0_n88_w70, c0_n88_w71, c0_n88_w72, c0_n88_w73, c0_n88_w74, c0_n88_w75, c0_n88_w76, c0_n88_w77, c0_n88_w78, c0_n88_w79, c0_n88_w80, c0_n88_w81, c0_n88_w82, c0_n88_w83, c0_n88_w84, c0_n88_w85, c0_n88_w86, c0_n88_w87, c0_n88_w88, c0_n88_w89, c0_n88_w90, c0_n88_w91, c0_n88_w92, c0_n88_w93, c0_n88_w94, c0_n88_w95, c0_n88_w96, c0_n88_w97, c0_n88_w98, c0_n88_w99, c0_n88_w100, c0_n88_w101, c0_n88_w102, c0_n88_w103, c0_n88_w104, c0_n88_w105, c0_n88_w106, c0_n88_w107, c0_n88_w108, c0_n88_w109, c0_n88_w110, c0_n88_w111, c0_n88_w112, c0_n88_w113, c0_n88_w114, c0_n88_w115, c0_n88_w116, c0_n88_w117, c0_n88_w118, c0_n88_w119, c0_n88_w120, c0_n88_w121, c0_n88_w122, c0_n88_w123, c0_n88_w124, c0_n88_w125, c0_n88_w126, c0_n88_w127, c0_n88_w128, c0_n88_w129, c0_n88_w130, c0_n88_w131, c0_n88_w132, c0_n88_w133, c0_n88_w134, c0_n88_w135, c0_n88_w136, c0_n88_w137, c0_n88_w138, c0_n88_w139, c0_n88_w140, c0_n88_w141, c0_n88_w142, c0_n88_w143, c0_n88_w144, c0_n88_w145, c0_n88_w146, c0_n88_w147, c0_n88_w148, c0_n88_w149, c0_n88_w150, c0_n88_w151, c0_n88_w152, c0_n88_w153, c0_n88_w154, c0_n88_w155, c0_n88_w156, c0_n88_w157, c0_n88_w158, c0_n88_w159, c0_n88_w160, c0_n88_w161, c0_n88_w162, c0_n88_w163, c0_n88_w164, c0_n88_w165, c0_n88_w166, c0_n88_w167, c0_n88_w168, c0_n88_w169, c0_n88_w170, c0_n88_w171, c0_n88_w172, c0_n88_w173, c0_n88_w174, c0_n88_w175, c0_n88_w176, c0_n88_w177, c0_n88_w178, c0_n88_w179, c0_n88_w180, c0_n88_w181, c0_n88_w182, c0_n88_w183, c0_n88_w184, c0_n88_w185, c0_n88_w186, c0_n88_w187, c0_n88_w188, c0_n88_w189, c0_n88_w190, c0_n88_w191, c0_n88_w192, c0_n88_w193, c0_n88_w194, c0_n88_w195, c0_n88_w196, c0_n88_w197, c0_n88_w198, c0_n88_w199, c0_n88_w200, c0_n89_w1, c0_n89_w2, c0_n89_w3, c0_n89_w4, c0_n89_w5, c0_n89_w6, c0_n89_w7, c0_n89_w8, c0_n89_w9, c0_n89_w10, c0_n89_w11, c0_n89_w12, c0_n89_w13, c0_n89_w14, c0_n89_w15, c0_n89_w16, c0_n89_w17, c0_n89_w18, c0_n89_w19, c0_n89_w20, c0_n89_w21, c0_n89_w22, c0_n89_w23, c0_n89_w24, c0_n89_w25, c0_n89_w26, c0_n89_w27, c0_n89_w28, c0_n89_w29, c0_n89_w30, c0_n89_w31, c0_n89_w32, c0_n89_w33, c0_n89_w34, c0_n89_w35, c0_n89_w36, c0_n89_w37, c0_n89_w38, c0_n89_w39, c0_n89_w40, c0_n89_w41, c0_n89_w42, c0_n89_w43, c0_n89_w44, c0_n89_w45, c0_n89_w46, c0_n89_w47, c0_n89_w48, c0_n89_w49, c0_n89_w50, c0_n89_w51, c0_n89_w52, c0_n89_w53, c0_n89_w54, c0_n89_w55, c0_n89_w56, c0_n89_w57, c0_n89_w58, c0_n89_w59, c0_n89_w60, c0_n89_w61, c0_n89_w62, c0_n89_w63, c0_n89_w64, c0_n89_w65, c0_n89_w66, c0_n89_w67, c0_n89_w68, c0_n89_w69, c0_n89_w70, c0_n89_w71, c0_n89_w72, c0_n89_w73, c0_n89_w74, c0_n89_w75, c0_n89_w76, c0_n89_w77, c0_n89_w78, c0_n89_w79, c0_n89_w80, c0_n89_w81, c0_n89_w82, c0_n89_w83, c0_n89_w84, c0_n89_w85, c0_n89_w86, c0_n89_w87, c0_n89_w88, c0_n89_w89, c0_n89_w90, c0_n89_w91, c0_n89_w92, c0_n89_w93, c0_n89_w94, c0_n89_w95, c0_n89_w96, c0_n89_w97, c0_n89_w98, c0_n89_w99, c0_n89_w100, c0_n89_w101, c0_n89_w102, c0_n89_w103, c0_n89_w104, c0_n89_w105, c0_n89_w106, c0_n89_w107, c0_n89_w108, c0_n89_w109, c0_n89_w110, c0_n89_w111, c0_n89_w112, c0_n89_w113, c0_n89_w114, c0_n89_w115, c0_n89_w116, c0_n89_w117, c0_n89_w118, c0_n89_w119, c0_n89_w120, c0_n89_w121, c0_n89_w122, c0_n89_w123, c0_n89_w124, c0_n89_w125, c0_n89_w126, c0_n89_w127, c0_n89_w128, c0_n89_w129, c0_n89_w130, c0_n89_w131, c0_n89_w132, c0_n89_w133, c0_n89_w134, c0_n89_w135, c0_n89_w136, c0_n89_w137, c0_n89_w138, c0_n89_w139, c0_n89_w140, c0_n89_w141, c0_n89_w142, c0_n89_w143, c0_n89_w144, c0_n89_w145, c0_n89_w146, c0_n89_w147, c0_n89_w148, c0_n89_w149, c0_n89_w150, c0_n89_w151, c0_n89_w152, c0_n89_w153, c0_n89_w154, c0_n89_w155, c0_n89_w156, c0_n89_w157, c0_n89_w158, c0_n89_w159, c0_n89_w160, c0_n89_w161, c0_n89_w162, c0_n89_w163, c0_n89_w164, c0_n89_w165, c0_n89_w166, c0_n89_w167, c0_n89_w168, c0_n89_w169, c0_n89_w170, c0_n89_w171, c0_n89_w172, c0_n89_w173, c0_n89_w174, c0_n89_w175, c0_n89_w176, c0_n89_w177, c0_n89_w178, c0_n89_w179, c0_n89_w180, c0_n89_w181, c0_n89_w182, c0_n89_w183, c0_n89_w184, c0_n89_w185, c0_n89_w186, c0_n89_w187, c0_n89_w188, c0_n89_w189, c0_n89_w190, c0_n89_w191, c0_n89_w192, c0_n89_w193, c0_n89_w194, c0_n89_w195, c0_n89_w196, c0_n89_w197, c0_n89_w198, c0_n89_w199, c0_n89_w200, c0_n90_w1, c0_n90_w2, c0_n90_w3, c0_n90_w4, c0_n90_w5, c0_n90_w6, c0_n90_w7, c0_n90_w8, c0_n90_w9, c0_n90_w10, c0_n90_w11, c0_n90_w12, c0_n90_w13, c0_n90_w14, c0_n90_w15, c0_n90_w16, c0_n90_w17, c0_n90_w18, c0_n90_w19, c0_n90_w20, c0_n90_w21, c0_n90_w22, c0_n90_w23, c0_n90_w24, c0_n90_w25, c0_n90_w26, c0_n90_w27, c0_n90_w28, c0_n90_w29, c0_n90_w30, c0_n90_w31, c0_n90_w32, c0_n90_w33, c0_n90_w34, c0_n90_w35, c0_n90_w36, c0_n90_w37, c0_n90_w38, c0_n90_w39, c0_n90_w40, c0_n90_w41, c0_n90_w42, c0_n90_w43, c0_n90_w44, c0_n90_w45, c0_n90_w46, c0_n90_w47, c0_n90_w48, c0_n90_w49, c0_n90_w50, c0_n90_w51, c0_n90_w52, c0_n90_w53, c0_n90_w54, c0_n90_w55, c0_n90_w56, c0_n90_w57, c0_n90_w58, c0_n90_w59, c0_n90_w60, c0_n90_w61, c0_n90_w62, c0_n90_w63, c0_n90_w64, c0_n90_w65, c0_n90_w66, c0_n90_w67, c0_n90_w68, c0_n90_w69, c0_n90_w70, c0_n90_w71, c0_n90_w72, c0_n90_w73, c0_n90_w74, c0_n90_w75, c0_n90_w76, c0_n90_w77, c0_n90_w78, c0_n90_w79, c0_n90_w80, c0_n90_w81, c0_n90_w82, c0_n90_w83, c0_n90_w84, c0_n90_w85, c0_n90_w86, c0_n90_w87, c0_n90_w88, c0_n90_w89, c0_n90_w90, c0_n90_w91, c0_n90_w92, c0_n90_w93, c0_n90_w94, c0_n90_w95, c0_n90_w96, c0_n90_w97, c0_n90_w98, c0_n90_w99, c0_n90_w100, c0_n90_w101, c0_n90_w102, c0_n90_w103, c0_n90_w104, c0_n90_w105, c0_n90_w106, c0_n90_w107, c0_n90_w108, c0_n90_w109, c0_n90_w110, c0_n90_w111, c0_n90_w112, c0_n90_w113, c0_n90_w114, c0_n90_w115, c0_n90_w116, c0_n90_w117, c0_n90_w118, c0_n90_w119, c0_n90_w120, c0_n90_w121, c0_n90_w122, c0_n90_w123, c0_n90_w124, c0_n90_w125, c0_n90_w126, c0_n90_w127, c0_n90_w128, c0_n90_w129, c0_n90_w130, c0_n90_w131, c0_n90_w132, c0_n90_w133, c0_n90_w134, c0_n90_w135, c0_n90_w136, c0_n90_w137, c0_n90_w138, c0_n90_w139, c0_n90_w140, c0_n90_w141, c0_n90_w142, c0_n90_w143, c0_n90_w144, c0_n90_w145, c0_n90_w146, c0_n90_w147, c0_n90_w148, c0_n90_w149, c0_n90_w150, c0_n90_w151, c0_n90_w152, c0_n90_w153, c0_n90_w154, c0_n90_w155, c0_n90_w156, c0_n90_w157, c0_n90_w158, c0_n90_w159, c0_n90_w160, c0_n90_w161, c0_n90_w162, c0_n90_w163, c0_n90_w164, c0_n90_w165, c0_n90_w166, c0_n90_w167, c0_n90_w168, c0_n90_w169, c0_n90_w170, c0_n90_w171, c0_n90_w172, c0_n90_w173, c0_n90_w174, c0_n90_w175, c0_n90_w176, c0_n90_w177, c0_n90_w178, c0_n90_w179, c0_n90_w180, c0_n90_w181, c0_n90_w182, c0_n90_w183, c0_n90_w184, c0_n90_w185, c0_n90_w186, c0_n90_w187, c0_n90_w188, c0_n90_w189, c0_n90_w190, c0_n90_w191, c0_n90_w192, c0_n90_w193, c0_n90_w194, c0_n90_w195, c0_n90_w196, c0_n90_w197, c0_n90_w198, c0_n90_w199, c0_n90_w200, c0_n91_w1, c0_n91_w2, c0_n91_w3, c0_n91_w4, c0_n91_w5, c0_n91_w6, c0_n91_w7, c0_n91_w8, c0_n91_w9, c0_n91_w10, c0_n91_w11, c0_n91_w12, c0_n91_w13, c0_n91_w14, c0_n91_w15, c0_n91_w16, c0_n91_w17, c0_n91_w18, c0_n91_w19, c0_n91_w20, c0_n91_w21, c0_n91_w22, c0_n91_w23, c0_n91_w24, c0_n91_w25, c0_n91_w26, c0_n91_w27, c0_n91_w28, c0_n91_w29, c0_n91_w30, c0_n91_w31, c0_n91_w32, c0_n91_w33, c0_n91_w34, c0_n91_w35, c0_n91_w36, c0_n91_w37, c0_n91_w38, c0_n91_w39, c0_n91_w40, c0_n91_w41, c0_n91_w42, c0_n91_w43, c0_n91_w44, c0_n91_w45, c0_n91_w46, c0_n91_w47, c0_n91_w48, c0_n91_w49, c0_n91_w50, c0_n91_w51, c0_n91_w52, c0_n91_w53, c0_n91_w54, c0_n91_w55, c0_n91_w56, c0_n91_w57, c0_n91_w58, c0_n91_w59, c0_n91_w60, c0_n91_w61, c0_n91_w62, c0_n91_w63, c0_n91_w64, c0_n91_w65, c0_n91_w66, c0_n91_w67, c0_n91_w68, c0_n91_w69, c0_n91_w70, c0_n91_w71, c0_n91_w72, c0_n91_w73, c0_n91_w74, c0_n91_w75, c0_n91_w76, c0_n91_w77, c0_n91_w78, c0_n91_w79, c0_n91_w80, c0_n91_w81, c0_n91_w82, c0_n91_w83, c0_n91_w84, c0_n91_w85, c0_n91_w86, c0_n91_w87, c0_n91_w88, c0_n91_w89, c0_n91_w90, c0_n91_w91, c0_n91_w92, c0_n91_w93, c0_n91_w94, c0_n91_w95, c0_n91_w96, c0_n91_w97, c0_n91_w98, c0_n91_w99, c0_n91_w100, c0_n91_w101, c0_n91_w102, c0_n91_w103, c0_n91_w104, c0_n91_w105, c0_n91_w106, c0_n91_w107, c0_n91_w108, c0_n91_w109, c0_n91_w110, c0_n91_w111, c0_n91_w112, c0_n91_w113, c0_n91_w114, c0_n91_w115, c0_n91_w116, c0_n91_w117, c0_n91_w118, c0_n91_w119, c0_n91_w120, c0_n91_w121, c0_n91_w122, c0_n91_w123, c0_n91_w124, c0_n91_w125, c0_n91_w126, c0_n91_w127, c0_n91_w128, c0_n91_w129, c0_n91_w130, c0_n91_w131, c0_n91_w132, c0_n91_w133, c0_n91_w134, c0_n91_w135, c0_n91_w136, c0_n91_w137, c0_n91_w138, c0_n91_w139, c0_n91_w140, c0_n91_w141, c0_n91_w142, c0_n91_w143, c0_n91_w144, c0_n91_w145, c0_n91_w146, c0_n91_w147, c0_n91_w148, c0_n91_w149, c0_n91_w150, c0_n91_w151, c0_n91_w152, c0_n91_w153, c0_n91_w154, c0_n91_w155, c0_n91_w156, c0_n91_w157, c0_n91_w158, c0_n91_w159, c0_n91_w160, c0_n91_w161, c0_n91_w162, c0_n91_w163, c0_n91_w164, c0_n91_w165, c0_n91_w166, c0_n91_w167, c0_n91_w168, c0_n91_w169, c0_n91_w170, c0_n91_w171, c0_n91_w172, c0_n91_w173, c0_n91_w174, c0_n91_w175, c0_n91_w176, c0_n91_w177, c0_n91_w178, c0_n91_w179, c0_n91_w180, c0_n91_w181, c0_n91_w182, c0_n91_w183, c0_n91_w184, c0_n91_w185, c0_n91_w186, c0_n91_w187, c0_n91_w188, c0_n91_w189, c0_n91_w190, c0_n91_w191, c0_n91_w192, c0_n91_w193, c0_n91_w194, c0_n91_w195, c0_n91_w196, c0_n91_w197, c0_n91_w198, c0_n91_w199, c0_n91_w200, c0_n92_w1, c0_n92_w2, c0_n92_w3, c0_n92_w4, c0_n92_w5, c0_n92_w6, c0_n92_w7, c0_n92_w8, c0_n92_w9, c0_n92_w10, c0_n92_w11, c0_n92_w12, c0_n92_w13, c0_n92_w14, c0_n92_w15, c0_n92_w16, c0_n92_w17, c0_n92_w18, c0_n92_w19, c0_n92_w20, c0_n92_w21, c0_n92_w22, c0_n92_w23, c0_n92_w24, c0_n92_w25, c0_n92_w26, c0_n92_w27, c0_n92_w28, c0_n92_w29, c0_n92_w30, c0_n92_w31, c0_n92_w32, c0_n92_w33, c0_n92_w34, c0_n92_w35, c0_n92_w36, c0_n92_w37, c0_n92_w38, c0_n92_w39, c0_n92_w40, c0_n92_w41, c0_n92_w42, c0_n92_w43, c0_n92_w44, c0_n92_w45, c0_n92_w46, c0_n92_w47, c0_n92_w48, c0_n92_w49, c0_n92_w50, c0_n92_w51, c0_n92_w52, c0_n92_w53, c0_n92_w54, c0_n92_w55, c0_n92_w56, c0_n92_w57, c0_n92_w58, c0_n92_w59, c0_n92_w60, c0_n92_w61, c0_n92_w62, c0_n92_w63, c0_n92_w64, c0_n92_w65, c0_n92_w66, c0_n92_w67, c0_n92_w68, c0_n92_w69, c0_n92_w70, c0_n92_w71, c0_n92_w72, c0_n92_w73, c0_n92_w74, c0_n92_w75, c0_n92_w76, c0_n92_w77, c0_n92_w78, c0_n92_w79, c0_n92_w80, c0_n92_w81, c0_n92_w82, c0_n92_w83, c0_n92_w84, c0_n92_w85, c0_n92_w86, c0_n92_w87, c0_n92_w88, c0_n92_w89, c0_n92_w90, c0_n92_w91, c0_n92_w92, c0_n92_w93, c0_n92_w94, c0_n92_w95, c0_n92_w96, c0_n92_w97, c0_n92_w98, c0_n92_w99, c0_n92_w100, c0_n92_w101, c0_n92_w102, c0_n92_w103, c0_n92_w104, c0_n92_w105, c0_n92_w106, c0_n92_w107, c0_n92_w108, c0_n92_w109, c0_n92_w110, c0_n92_w111, c0_n92_w112, c0_n92_w113, c0_n92_w114, c0_n92_w115, c0_n92_w116, c0_n92_w117, c0_n92_w118, c0_n92_w119, c0_n92_w120, c0_n92_w121, c0_n92_w122, c0_n92_w123, c0_n92_w124, c0_n92_w125, c0_n92_w126, c0_n92_w127, c0_n92_w128, c0_n92_w129, c0_n92_w130, c0_n92_w131, c0_n92_w132, c0_n92_w133, c0_n92_w134, c0_n92_w135, c0_n92_w136, c0_n92_w137, c0_n92_w138, c0_n92_w139, c0_n92_w140, c0_n92_w141, c0_n92_w142, c0_n92_w143, c0_n92_w144, c0_n92_w145, c0_n92_w146, c0_n92_w147, c0_n92_w148, c0_n92_w149, c0_n92_w150, c0_n92_w151, c0_n92_w152, c0_n92_w153, c0_n92_w154, c0_n92_w155, c0_n92_w156, c0_n92_w157, c0_n92_w158, c0_n92_w159, c0_n92_w160, c0_n92_w161, c0_n92_w162, c0_n92_w163, c0_n92_w164, c0_n92_w165, c0_n92_w166, c0_n92_w167, c0_n92_w168, c0_n92_w169, c0_n92_w170, c0_n92_w171, c0_n92_w172, c0_n92_w173, c0_n92_w174, c0_n92_w175, c0_n92_w176, c0_n92_w177, c0_n92_w178, c0_n92_w179, c0_n92_w180, c0_n92_w181, c0_n92_w182, c0_n92_w183, c0_n92_w184, c0_n92_w185, c0_n92_w186, c0_n92_w187, c0_n92_w188, c0_n92_w189, c0_n92_w190, c0_n92_w191, c0_n92_w192, c0_n92_w193, c0_n92_w194, c0_n92_w195, c0_n92_w196, c0_n92_w197, c0_n92_w198, c0_n92_w199, c0_n92_w200, c0_n93_w1, c0_n93_w2, c0_n93_w3, c0_n93_w4, c0_n93_w5, c0_n93_w6, c0_n93_w7, c0_n93_w8, c0_n93_w9, c0_n93_w10, c0_n93_w11, c0_n93_w12, c0_n93_w13, c0_n93_w14, c0_n93_w15, c0_n93_w16, c0_n93_w17, c0_n93_w18, c0_n93_w19, c0_n93_w20, c0_n93_w21, c0_n93_w22, c0_n93_w23, c0_n93_w24, c0_n93_w25, c0_n93_w26, c0_n93_w27, c0_n93_w28, c0_n93_w29, c0_n93_w30, c0_n93_w31, c0_n93_w32, c0_n93_w33, c0_n93_w34, c0_n93_w35, c0_n93_w36, c0_n93_w37, c0_n93_w38, c0_n93_w39, c0_n93_w40, c0_n93_w41, c0_n93_w42, c0_n93_w43, c0_n93_w44, c0_n93_w45, c0_n93_w46, c0_n93_w47, c0_n93_w48, c0_n93_w49, c0_n93_w50, c0_n93_w51, c0_n93_w52, c0_n93_w53, c0_n93_w54, c0_n93_w55, c0_n93_w56, c0_n93_w57, c0_n93_w58, c0_n93_w59, c0_n93_w60, c0_n93_w61, c0_n93_w62, c0_n93_w63, c0_n93_w64, c0_n93_w65, c0_n93_w66, c0_n93_w67, c0_n93_w68, c0_n93_w69, c0_n93_w70, c0_n93_w71, c0_n93_w72, c0_n93_w73, c0_n93_w74, c0_n93_w75, c0_n93_w76, c0_n93_w77, c0_n93_w78, c0_n93_w79, c0_n93_w80, c0_n93_w81, c0_n93_w82, c0_n93_w83, c0_n93_w84, c0_n93_w85, c0_n93_w86, c0_n93_w87, c0_n93_w88, c0_n93_w89, c0_n93_w90, c0_n93_w91, c0_n93_w92, c0_n93_w93, c0_n93_w94, c0_n93_w95, c0_n93_w96, c0_n93_w97, c0_n93_w98, c0_n93_w99, c0_n93_w100, c0_n93_w101, c0_n93_w102, c0_n93_w103, c0_n93_w104, c0_n93_w105, c0_n93_w106, c0_n93_w107, c0_n93_w108, c0_n93_w109, c0_n93_w110, c0_n93_w111, c0_n93_w112, c0_n93_w113, c0_n93_w114, c0_n93_w115, c0_n93_w116, c0_n93_w117, c0_n93_w118, c0_n93_w119, c0_n93_w120, c0_n93_w121, c0_n93_w122, c0_n93_w123, c0_n93_w124, c0_n93_w125, c0_n93_w126, c0_n93_w127, c0_n93_w128, c0_n93_w129, c0_n93_w130, c0_n93_w131, c0_n93_w132, c0_n93_w133, c0_n93_w134, c0_n93_w135, c0_n93_w136, c0_n93_w137, c0_n93_w138, c0_n93_w139, c0_n93_w140, c0_n93_w141, c0_n93_w142, c0_n93_w143, c0_n93_w144, c0_n93_w145, c0_n93_w146, c0_n93_w147, c0_n93_w148, c0_n93_w149, c0_n93_w150, c0_n93_w151, c0_n93_w152, c0_n93_w153, c0_n93_w154, c0_n93_w155, c0_n93_w156, c0_n93_w157, c0_n93_w158, c0_n93_w159, c0_n93_w160, c0_n93_w161, c0_n93_w162, c0_n93_w163, c0_n93_w164, c0_n93_w165, c0_n93_w166, c0_n93_w167, c0_n93_w168, c0_n93_w169, c0_n93_w170, c0_n93_w171, c0_n93_w172, c0_n93_w173, c0_n93_w174, c0_n93_w175, c0_n93_w176, c0_n93_w177, c0_n93_w178, c0_n93_w179, c0_n93_w180, c0_n93_w181, c0_n93_w182, c0_n93_w183, c0_n93_w184, c0_n93_w185, c0_n93_w186, c0_n93_w187, c0_n93_w188, c0_n93_w189, c0_n93_w190, c0_n93_w191, c0_n93_w192, c0_n93_w193, c0_n93_w194, c0_n93_w195, c0_n93_w196, c0_n93_w197, c0_n93_w198, c0_n93_w199, c0_n93_w200, c0_n94_w1, c0_n94_w2, c0_n94_w3, c0_n94_w4, c0_n94_w5, c0_n94_w6, c0_n94_w7, c0_n94_w8, c0_n94_w9, c0_n94_w10, c0_n94_w11, c0_n94_w12, c0_n94_w13, c0_n94_w14, c0_n94_w15, c0_n94_w16, c0_n94_w17, c0_n94_w18, c0_n94_w19, c0_n94_w20, c0_n94_w21, c0_n94_w22, c0_n94_w23, c0_n94_w24, c0_n94_w25, c0_n94_w26, c0_n94_w27, c0_n94_w28, c0_n94_w29, c0_n94_w30, c0_n94_w31, c0_n94_w32, c0_n94_w33, c0_n94_w34, c0_n94_w35, c0_n94_w36, c0_n94_w37, c0_n94_w38, c0_n94_w39, c0_n94_w40, c0_n94_w41, c0_n94_w42, c0_n94_w43, c0_n94_w44, c0_n94_w45, c0_n94_w46, c0_n94_w47, c0_n94_w48, c0_n94_w49, c0_n94_w50, c0_n94_w51, c0_n94_w52, c0_n94_w53, c0_n94_w54, c0_n94_w55, c0_n94_w56, c0_n94_w57, c0_n94_w58, c0_n94_w59, c0_n94_w60, c0_n94_w61, c0_n94_w62, c0_n94_w63, c0_n94_w64, c0_n94_w65, c0_n94_w66, c0_n94_w67, c0_n94_w68, c0_n94_w69, c0_n94_w70, c0_n94_w71, c0_n94_w72, c0_n94_w73, c0_n94_w74, c0_n94_w75, c0_n94_w76, c0_n94_w77, c0_n94_w78, c0_n94_w79, c0_n94_w80, c0_n94_w81, c0_n94_w82, c0_n94_w83, c0_n94_w84, c0_n94_w85, c0_n94_w86, c0_n94_w87, c0_n94_w88, c0_n94_w89, c0_n94_w90, c0_n94_w91, c0_n94_w92, c0_n94_w93, c0_n94_w94, c0_n94_w95, c0_n94_w96, c0_n94_w97, c0_n94_w98, c0_n94_w99, c0_n94_w100, c0_n94_w101, c0_n94_w102, c0_n94_w103, c0_n94_w104, c0_n94_w105, c0_n94_w106, c0_n94_w107, c0_n94_w108, c0_n94_w109, c0_n94_w110, c0_n94_w111, c0_n94_w112, c0_n94_w113, c0_n94_w114, c0_n94_w115, c0_n94_w116, c0_n94_w117, c0_n94_w118, c0_n94_w119, c0_n94_w120, c0_n94_w121, c0_n94_w122, c0_n94_w123, c0_n94_w124, c0_n94_w125, c0_n94_w126, c0_n94_w127, c0_n94_w128, c0_n94_w129, c0_n94_w130, c0_n94_w131, c0_n94_w132, c0_n94_w133, c0_n94_w134, c0_n94_w135, c0_n94_w136, c0_n94_w137, c0_n94_w138, c0_n94_w139, c0_n94_w140, c0_n94_w141, c0_n94_w142, c0_n94_w143, c0_n94_w144, c0_n94_w145, c0_n94_w146, c0_n94_w147, c0_n94_w148, c0_n94_w149, c0_n94_w150, c0_n94_w151, c0_n94_w152, c0_n94_w153, c0_n94_w154, c0_n94_w155, c0_n94_w156, c0_n94_w157, c0_n94_w158, c0_n94_w159, c0_n94_w160, c0_n94_w161, c0_n94_w162, c0_n94_w163, c0_n94_w164, c0_n94_w165, c0_n94_w166, c0_n94_w167, c0_n94_w168, c0_n94_w169, c0_n94_w170, c0_n94_w171, c0_n94_w172, c0_n94_w173, c0_n94_w174, c0_n94_w175, c0_n94_w176, c0_n94_w177, c0_n94_w178, c0_n94_w179, c0_n94_w180, c0_n94_w181, c0_n94_w182, c0_n94_w183, c0_n94_w184, c0_n94_w185, c0_n94_w186, c0_n94_w187, c0_n94_w188, c0_n94_w189, c0_n94_w190, c0_n94_w191, c0_n94_w192, c0_n94_w193, c0_n94_w194, c0_n94_w195, c0_n94_w196, c0_n94_w197, c0_n94_w198, c0_n94_w199, c0_n94_w200, c0_n95_w1, c0_n95_w2, c0_n95_w3, c0_n95_w4, c0_n95_w5, c0_n95_w6, c0_n95_w7, c0_n95_w8, c0_n95_w9, c0_n95_w10, c0_n95_w11, c0_n95_w12, c0_n95_w13, c0_n95_w14, c0_n95_w15, c0_n95_w16, c0_n95_w17, c0_n95_w18, c0_n95_w19, c0_n95_w20, c0_n95_w21, c0_n95_w22, c0_n95_w23, c0_n95_w24, c0_n95_w25, c0_n95_w26, c0_n95_w27, c0_n95_w28, c0_n95_w29, c0_n95_w30, c0_n95_w31, c0_n95_w32, c0_n95_w33, c0_n95_w34, c0_n95_w35, c0_n95_w36, c0_n95_w37, c0_n95_w38, c0_n95_w39, c0_n95_w40, c0_n95_w41, c0_n95_w42, c0_n95_w43, c0_n95_w44, c0_n95_w45, c0_n95_w46, c0_n95_w47, c0_n95_w48, c0_n95_w49, c0_n95_w50, c0_n95_w51, c0_n95_w52, c0_n95_w53, c0_n95_w54, c0_n95_w55, c0_n95_w56, c0_n95_w57, c0_n95_w58, c0_n95_w59, c0_n95_w60, c0_n95_w61, c0_n95_w62, c0_n95_w63, c0_n95_w64, c0_n95_w65, c0_n95_w66, c0_n95_w67, c0_n95_w68, c0_n95_w69, c0_n95_w70, c0_n95_w71, c0_n95_w72, c0_n95_w73, c0_n95_w74, c0_n95_w75, c0_n95_w76, c0_n95_w77, c0_n95_w78, c0_n95_w79, c0_n95_w80, c0_n95_w81, c0_n95_w82, c0_n95_w83, c0_n95_w84, c0_n95_w85, c0_n95_w86, c0_n95_w87, c0_n95_w88, c0_n95_w89, c0_n95_w90, c0_n95_w91, c0_n95_w92, c0_n95_w93, c0_n95_w94, c0_n95_w95, c0_n95_w96, c0_n95_w97, c0_n95_w98, c0_n95_w99, c0_n95_w100, c0_n95_w101, c0_n95_w102, c0_n95_w103, c0_n95_w104, c0_n95_w105, c0_n95_w106, c0_n95_w107, c0_n95_w108, c0_n95_w109, c0_n95_w110, c0_n95_w111, c0_n95_w112, c0_n95_w113, c0_n95_w114, c0_n95_w115, c0_n95_w116, c0_n95_w117, c0_n95_w118, c0_n95_w119, c0_n95_w120, c0_n95_w121, c0_n95_w122, c0_n95_w123, c0_n95_w124, c0_n95_w125, c0_n95_w126, c0_n95_w127, c0_n95_w128, c0_n95_w129, c0_n95_w130, c0_n95_w131, c0_n95_w132, c0_n95_w133, c0_n95_w134, c0_n95_w135, c0_n95_w136, c0_n95_w137, c0_n95_w138, c0_n95_w139, c0_n95_w140, c0_n95_w141, c0_n95_w142, c0_n95_w143, c0_n95_w144, c0_n95_w145, c0_n95_w146, c0_n95_w147, c0_n95_w148, c0_n95_w149, c0_n95_w150, c0_n95_w151, c0_n95_w152, c0_n95_w153, c0_n95_w154, c0_n95_w155, c0_n95_w156, c0_n95_w157, c0_n95_w158, c0_n95_w159, c0_n95_w160, c0_n95_w161, c0_n95_w162, c0_n95_w163, c0_n95_w164, c0_n95_w165, c0_n95_w166, c0_n95_w167, c0_n95_w168, c0_n95_w169, c0_n95_w170, c0_n95_w171, c0_n95_w172, c0_n95_w173, c0_n95_w174, c0_n95_w175, c0_n95_w176, c0_n95_w177, c0_n95_w178, c0_n95_w179, c0_n95_w180, c0_n95_w181, c0_n95_w182, c0_n95_w183, c0_n95_w184, c0_n95_w185, c0_n95_w186, c0_n95_w187, c0_n95_w188, c0_n95_w189, c0_n95_w190, c0_n95_w191, c0_n95_w192, c0_n95_w193, c0_n95_w194, c0_n95_w195, c0_n95_w196, c0_n95_w197, c0_n95_w198, c0_n95_w199, c0_n95_w200, c0_n96_w1, c0_n96_w2, c0_n96_w3, c0_n96_w4, c0_n96_w5, c0_n96_w6, c0_n96_w7, c0_n96_w8, c0_n96_w9, c0_n96_w10, c0_n96_w11, c0_n96_w12, c0_n96_w13, c0_n96_w14, c0_n96_w15, c0_n96_w16, c0_n96_w17, c0_n96_w18, c0_n96_w19, c0_n96_w20, c0_n96_w21, c0_n96_w22, c0_n96_w23, c0_n96_w24, c0_n96_w25, c0_n96_w26, c0_n96_w27, c0_n96_w28, c0_n96_w29, c0_n96_w30, c0_n96_w31, c0_n96_w32, c0_n96_w33, c0_n96_w34, c0_n96_w35, c0_n96_w36, c0_n96_w37, c0_n96_w38, c0_n96_w39, c0_n96_w40, c0_n96_w41, c0_n96_w42, c0_n96_w43, c0_n96_w44, c0_n96_w45, c0_n96_w46, c0_n96_w47, c0_n96_w48, c0_n96_w49, c0_n96_w50, c0_n96_w51, c0_n96_w52, c0_n96_w53, c0_n96_w54, c0_n96_w55, c0_n96_w56, c0_n96_w57, c0_n96_w58, c0_n96_w59, c0_n96_w60, c0_n96_w61, c0_n96_w62, c0_n96_w63, c0_n96_w64, c0_n96_w65, c0_n96_w66, c0_n96_w67, c0_n96_w68, c0_n96_w69, c0_n96_w70, c0_n96_w71, c0_n96_w72, c0_n96_w73, c0_n96_w74, c0_n96_w75, c0_n96_w76, c0_n96_w77, c0_n96_w78, c0_n96_w79, c0_n96_w80, c0_n96_w81, c0_n96_w82, c0_n96_w83, c0_n96_w84, c0_n96_w85, c0_n96_w86, c0_n96_w87, c0_n96_w88, c0_n96_w89, c0_n96_w90, c0_n96_w91, c0_n96_w92, c0_n96_w93, c0_n96_w94, c0_n96_w95, c0_n96_w96, c0_n96_w97, c0_n96_w98, c0_n96_w99, c0_n96_w100, c0_n96_w101, c0_n96_w102, c0_n96_w103, c0_n96_w104, c0_n96_w105, c0_n96_w106, c0_n96_w107, c0_n96_w108, c0_n96_w109, c0_n96_w110, c0_n96_w111, c0_n96_w112, c0_n96_w113, c0_n96_w114, c0_n96_w115, c0_n96_w116, c0_n96_w117, c0_n96_w118, c0_n96_w119, c0_n96_w120, c0_n96_w121, c0_n96_w122, c0_n96_w123, c0_n96_w124, c0_n96_w125, c0_n96_w126, c0_n96_w127, c0_n96_w128, c0_n96_w129, c0_n96_w130, c0_n96_w131, c0_n96_w132, c0_n96_w133, c0_n96_w134, c0_n96_w135, c0_n96_w136, c0_n96_w137, c0_n96_w138, c0_n96_w139, c0_n96_w140, c0_n96_w141, c0_n96_w142, c0_n96_w143, c0_n96_w144, c0_n96_w145, c0_n96_w146, c0_n96_w147, c0_n96_w148, c0_n96_w149, c0_n96_w150, c0_n96_w151, c0_n96_w152, c0_n96_w153, c0_n96_w154, c0_n96_w155, c0_n96_w156, c0_n96_w157, c0_n96_w158, c0_n96_w159, c0_n96_w160, c0_n96_w161, c0_n96_w162, c0_n96_w163, c0_n96_w164, c0_n96_w165, c0_n96_w166, c0_n96_w167, c0_n96_w168, c0_n96_w169, c0_n96_w170, c0_n96_w171, c0_n96_w172, c0_n96_w173, c0_n96_w174, c0_n96_w175, c0_n96_w176, c0_n96_w177, c0_n96_w178, c0_n96_w179, c0_n96_w180, c0_n96_w181, c0_n96_w182, c0_n96_w183, c0_n96_w184, c0_n96_w185, c0_n96_w186, c0_n96_w187, c0_n96_w188, c0_n96_w189, c0_n96_w190, c0_n96_w191, c0_n96_w192, c0_n96_w193, c0_n96_w194, c0_n96_w195, c0_n96_w196, c0_n96_w197, c0_n96_w198, c0_n96_w199, c0_n96_w200, c0_n97_w1, c0_n97_w2, c0_n97_w3, c0_n97_w4, c0_n97_w5, c0_n97_w6, c0_n97_w7, c0_n97_w8, c0_n97_w9, c0_n97_w10, c0_n97_w11, c0_n97_w12, c0_n97_w13, c0_n97_w14, c0_n97_w15, c0_n97_w16, c0_n97_w17, c0_n97_w18, c0_n97_w19, c0_n97_w20, c0_n97_w21, c0_n97_w22, c0_n97_w23, c0_n97_w24, c0_n97_w25, c0_n97_w26, c0_n97_w27, c0_n97_w28, c0_n97_w29, c0_n97_w30, c0_n97_w31, c0_n97_w32, c0_n97_w33, c0_n97_w34, c0_n97_w35, c0_n97_w36, c0_n97_w37, c0_n97_w38, c0_n97_w39, c0_n97_w40, c0_n97_w41, c0_n97_w42, c0_n97_w43, c0_n97_w44, c0_n97_w45, c0_n97_w46, c0_n97_w47, c0_n97_w48, c0_n97_w49, c0_n97_w50, c0_n97_w51, c0_n97_w52, c0_n97_w53, c0_n97_w54, c0_n97_w55, c0_n97_w56, c0_n97_w57, c0_n97_w58, c0_n97_w59, c0_n97_w60, c0_n97_w61, c0_n97_w62, c0_n97_w63, c0_n97_w64, c0_n97_w65, c0_n97_w66, c0_n97_w67, c0_n97_w68, c0_n97_w69, c0_n97_w70, c0_n97_w71, c0_n97_w72, c0_n97_w73, c0_n97_w74, c0_n97_w75, c0_n97_w76, c0_n97_w77, c0_n97_w78, c0_n97_w79, c0_n97_w80, c0_n97_w81, c0_n97_w82, c0_n97_w83, c0_n97_w84, c0_n97_w85, c0_n97_w86, c0_n97_w87, c0_n97_w88, c0_n97_w89, c0_n97_w90, c0_n97_w91, c0_n97_w92, c0_n97_w93, c0_n97_w94, c0_n97_w95, c0_n97_w96, c0_n97_w97, c0_n97_w98, c0_n97_w99, c0_n97_w100, c0_n97_w101, c0_n97_w102, c0_n97_w103, c0_n97_w104, c0_n97_w105, c0_n97_w106, c0_n97_w107, c0_n97_w108, c0_n97_w109, c0_n97_w110, c0_n97_w111, c0_n97_w112, c0_n97_w113, c0_n97_w114, c0_n97_w115, c0_n97_w116, c0_n97_w117, c0_n97_w118, c0_n97_w119, c0_n97_w120, c0_n97_w121, c0_n97_w122, c0_n97_w123, c0_n97_w124, c0_n97_w125, c0_n97_w126, c0_n97_w127, c0_n97_w128, c0_n97_w129, c0_n97_w130, c0_n97_w131, c0_n97_w132, c0_n97_w133, c0_n97_w134, c0_n97_w135, c0_n97_w136, c0_n97_w137, c0_n97_w138, c0_n97_w139, c0_n97_w140, c0_n97_w141, c0_n97_w142, c0_n97_w143, c0_n97_w144, c0_n97_w145, c0_n97_w146, c0_n97_w147, c0_n97_w148, c0_n97_w149, c0_n97_w150, c0_n97_w151, c0_n97_w152, c0_n97_w153, c0_n97_w154, c0_n97_w155, c0_n97_w156, c0_n97_w157, c0_n97_w158, c0_n97_w159, c0_n97_w160, c0_n97_w161, c0_n97_w162, c0_n97_w163, c0_n97_w164, c0_n97_w165, c0_n97_w166, c0_n97_w167, c0_n97_w168, c0_n97_w169, c0_n97_w170, c0_n97_w171, c0_n97_w172, c0_n97_w173, c0_n97_w174, c0_n97_w175, c0_n97_w176, c0_n97_w177, c0_n97_w178, c0_n97_w179, c0_n97_w180, c0_n97_w181, c0_n97_w182, c0_n97_w183, c0_n97_w184, c0_n97_w185, c0_n97_w186, c0_n97_w187, c0_n97_w188, c0_n97_w189, c0_n97_w190, c0_n97_w191, c0_n97_w192, c0_n97_w193, c0_n97_w194, c0_n97_w195, c0_n97_w196, c0_n97_w197, c0_n97_w198, c0_n97_w199, c0_n97_w200, c0_n98_w1, c0_n98_w2, c0_n98_w3, c0_n98_w4, c0_n98_w5, c0_n98_w6, c0_n98_w7, c0_n98_w8, c0_n98_w9, c0_n98_w10, c0_n98_w11, c0_n98_w12, c0_n98_w13, c0_n98_w14, c0_n98_w15, c0_n98_w16, c0_n98_w17, c0_n98_w18, c0_n98_w19, c0_n98_w20, c0_n98_w21, c0_n98_w22, c0_n98_w23, c0_n98_w24, c0_n98_w25, c0_n98_w26, c0_n98_w27, c0_n98_w28, c0_n98_w29, c0_n98_w30, c0_n98_w31, c0_n98_w32, c0_n98_w33, c0_n98_w34, c0_n98_w35, c0_n98_w36, c0_n98_w37, c0_n98_w38, c0_n98_w39, c0_n98_w40, c0_n98_w41, c0_n98_w42, c0_n98_w43, c0_n98_w44, c0_n98_w45, c0_n98_w46, c0_n98_w47, c0_n98_w48, c0_n98_w49, c0_n98_w50, c0_n98_w51, c0_n98_w52, c0_n98_w53, c0_n98_w54, c0_n98_w55, c0_n98_w56, c0_n98_w57, c0_n98_w58, c0_n98_w59, c0_n98_w60, c0_n98_w61, c0_n98_w62, c0_n98_w63, c0_n98_w64, c0_n98_w65, c0_n98_w66, c0_n98_w67, c0_n98_w68, c0_n98_w69, c0_n98_w70, c0_n98_w71, c0_n98_w72, c0_n98_w73, c0_n98_w74, c0_n98_w75, c0_n98_w76, c0_n98_w77, c0_n98_w78, c0_n98_w79, c0_n98_w80, c0_n98_w81, c0_n98_w82, c0_n98_w83, c0_n98_w84, c0_n98_w85, c0_n98_w86, c0_n98_w87, c0_n98_w88, c0_n98_w89, c0_n98_w90, c0_n98_w91, c0_n98_w92, c0_n98_w93, c0_n98_w94, c0_n98_w95, c0_n98_w96, c0_n98_w97, c0_n98_w98, c0_n98_w99, c0_n98_w100, c0_n98_w101, c0_n98_w102, c0_n98_w103, c0_n98_w104, c0_n98_w105, c0_n98_w106, c0_n98_w107, c0_n98_w108, c0_n98_w109, c0_n98_w110, c0_n98_w111, c0_n98_w112, c0_n98_w113, c0_n98_w114, c0_n98_w115, c0_n98_w116, c0_n98_w117, c0_n98_w118, c0_n98_w119, c0_n98_w120, c0_n98_w121, c0_n98_w122, c0_n98_w123, c0_n98_w124, c0_n98_w125, c0_n98_w126, c0_n98_w127, c0_n98_w128, c0_n98_w129, c0_n98_w130, c0_n98_w131, c0_n98_w132, c0_n98_w133, c0_n98_w134, c0_n98_w135, c0_n98_w136, c0_n98_w137, c0_n98_w138, c0_n98_w139, c0_n98_w140, c0_n98_w141, c0_n98_w142, c0_n98_w143, c0_n98_w144, c0_n98_w145, c0_n98_w146, c0_n98_w147, c0_n98_w148, c0_n98_w149, c0_n98_w150, c0_n98_w151, c0_n98_w152, c0_n98_w153, c0_n98_w154, c0_n98_w155, c0_n98_w156, c0_n98_w157, c0_n98_w158, c0_n98_w159, c0_n98_w160, c0_n98_w161, c0_n98_w162, c0_n98_w163, c0_n98_w164, c0_n98_w165, c0_n98_w166, c0_n98_w167, c0_n98_w168, c0_n98_w169, c0_n98_w170, c0_n98_w171, c0_n98_w172, c0_n98_w173, c0_n98_w174, c0_n98_w175, c0_n98_w176, c0_n98_w177, c0_n98_w178, c0_n98_w179, c0_n98_w180, c0_n98_w181, c0_n98_w182, c0_n98_w183, c0_n98_w184, c0_n98_w185, c0_n98_w186, c0_n98_w187, c0_n98_w188, c0_n98_w189, c0_n98_w190, c0_n98_w191, c0_n98_w192, c0_n98_w193, c0_n98_w194, c0_n98_w195, c0_n98_w196, c0_n98_w197, c0_n98_w198, c0_n98_w199, c0_n98_w200, c0_n99_w1, c0_n99_w2, c0_n99_w3, c0_n99_w4, c0_n99_w5, c0_n99_w6, c0_n99_w7, c0_n99_w8, c0_n99_w9, c0_n99_w10, c0_n99_w11, c0_n99_w12, c0_n99_w13, c0_n99_w14, c0_n99_w15, c0_n99_w16, c0_n99_w17, c0_n99_w18, c0_n99_w19, c0_n99_w20, c0_n99_w21, c0_n99_w22, c0_n99_w23, c0_n99_w24, c0_n99_w25, c0_n99_w26, c0_n99_w27, c0_n99_w28, c0_n99_w29, c0_n99_w30, c0_n99_w31, c0_n99_w32, c0_n99_w33, c0_n99_w34, c0_n99_w35, c0_n99_w36, c0_n99_w37, c0_n99_w38, c0_n99_w39, c0_n99_w40, c0_n99_w41, c0_n99_w42, c0_n99_w43, c0_n99_w44, c0_n99_w45, c0_n99_w46, c0_n99_w47, c0_n99_w48, c0_n99_w49, c0_n99_w50, c0_n99_w51, c0_n99_w52, c0_n99_w53, c0_n99_w54, c0_n99_w55, c0_n99_w56, c0_n99_w57, c0_n99_w58, c0_n99_w59, c0_n99_w60, c0_n99_w61, c0_n99_w62, c0_n99_w63, c0_n99_w64, c0_n99_w65, c0_n99_w66, c0_n99_w67, c0_n99_w68, c0_n99_w69, c0_n99_w70, c0_n99_w71, c0_n99_w72, c0_n99_w73, c0_n99_w74, c0_n99_w75, c0_n99_w76, c0_n99_w77, c0_n99_w78, c0_n99_w79, c0_n99_w80, c0_n99_w81, c0_n99_w82, c0_n99_w83, c0_n99_w84, c0_n99_w85, c0_n99_w86, c0_n99_w87, c0_n99_w88, c0_n99_w89, c0_n99_w90, c0_n99_w91, c0_n99_w92, c0_n99_w93, c0_n99_w94, c0_n99_w95, c0_n99_w96, c0_n99_w97, c0_n99_w98, c0_n99_w99, c0_n99_w100, c0_n99_w101, c0_n99_w102, c0_n99_w103, c0_n99_w104, c0_n99_w105, c0_n99_w106, c0_n99_w107, c0_n99_w108, c0_n99_w109, c0_n99_w110, c0_n99_w111, c0_n99_w112, c0_n99_w113, c0_n99_w114, c0_n99_w115, c0_n99_w116, c0_n99_w117, c0_n99_w118, c0_n99_w119, c0_n99_w120, c0_n99_w121, c0_n99_w122, c0_n99_w123, c0_n99_w124, c0_n99_w125, c0_n99_w126, c0_n99_w127, c0_n99_w128, c0_n99_w129, c0_n99_w130, c0_n99_w131, c0_n99_w132, c0_n99_w133, c0_n99_w134, c0_n99_w135, c0_n99_w136, c0_n99_w137, c0_n99_w138, c0_n99_w139, c0_n99_w140, c0_n99_w141, c0_n99_w142, c0_n99_w143, c0_n99_w144, c0_n99_w145, c0_n99_w146, c0_n99_w147, c0_n99_w148, c0_n99_w149, c0_n99_w150, c0_n99_w151, c0_n99_w152, c0_n99_w153, c0_n99_w154, c0_n99_w155, c0_n99_w156, c0_n99_w157, c0_n99_w158, c0_n99_w159, c0_n99_w160, c0_n99_w161, c0_n99_w162, c0_n99_w163, c0_n99_w164, c0_n99_w165, c0_n99_w166, c0_n99_w167, c0_n99_w168, c0_n99_w169, c0_n99_w170, c0_n99_w171, c0_n99_w172, c0_n99_w173, c0_n99_w174, c0_n99_w175, c0_n99_w176, c0_n99_w177, c0_n99_w178, c0_n99_w179, c0_n99_w180, c0_n99_w181, c0_n99_w182, c0_n99_w183, c0_n99_w184, c0_n99_w185, c0_n99_w186, c0_n99_w187, c0_n99_w188, c0_n99_w189, c0_n99_w190, c0_n99_w191, c0_n99_w192, c0_n99_w193, c0_n99_w194, c0_n99_w195, c0_n99_w196, c0_n99_w197, c0_n99_w198, c0_n99_w199, c0_n99_w200: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c0_n0_y, c0_n1_y, c0_n2_y, c0_n3_y, c0_n4_y, c0_n5_y, c0_n6_y, c0_n7_y, c0_n8_y, c0_n9_y, c0_n10_y, c0_n11_y, c0_n12_y, c0_n13_y, c0_n14_y, c0_n15_y, c0_n16_y, c0_n17_y, c0_n18_y, c0_n19_y, c0_n20_y, c0_n21_y, c0_n22_y, c0_n23_y, c0_n24_y, c0_n25_y, c0_n26_y, c0_n27_y, c0_n28_y, c0_n29_y, c0_n30_y, c0_n31_y, c0_n32_y, c0_n33_y, c0_n34_y, c0_n35_y, c0_n36_y, c0_n37_y, c0_n38_y, c0_n39_y, c0_n40_y, c0_n41_y, c0_n42_y, c0_n43_y, c0_n44_y, c0_n45_y, c0_n46_y, c0_n47_y, c0_n48_y, c0_n49_y, c0_n50_y, c0_n51_y, c0_n52_y, c0_n53_y, c0_n54_y, c0_n55_y, c0_n56_y, c0_n57_y, c0_n58_y, c0_n59_y, c0_n60_y, c0_n61_y, c0_n62_y, c0_n63_y, c0_n64_y, c0_n65_y, c0_n66_y, c0_n67_y, c0_n68_y, c0_n69_y, c0_n70_y, c0_n71_y, c0_n72_y, c0_n73_y, c0_n74_y, c0_n75_y, c0_n76_y, c0_n77_y, c0_n78_y, c0_n79_y, c0_n80_y, c0_n81_y, c0_n82_y, c0_n83_y, c0_n84_y, c0_n85_y, c0_n86_y, c0_n87_y, c0_n88_y, c0_n89_y, c0_n90_y, c0_n91_y, c0_n92_y, c0_n93_y, c0_n94_y, c0_n95_y, c0_n96_y, c0_n97_y, c0_n98_y, c0_n99_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada0_ReLU_100neuron_8bits_200n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n0_w1, 
            w2=> c0_n0_w2, 
            w3=> c0_n0_w3, 
            w4=> c0_n0_w4, 
            w5=> c0_n0_w5, 
            w6=> c0_n0_w6, 
            w7=> c0_n0_w7, 
            w8=> c0_n0_w8, 
            w9=> c0_n0_w9, 
            w10=> c0_n0_w10, 
            w11=> c0_n0_w11, 
            w12=> c0_n0_w12, 
            w13=> c0_n0_w13, 
            w14=> c0_n0_w14, 
            w15=> c0_n0_w15, 
            w16=> c0_n0_w16, 
            w17=> c0_n0_w17, 
            w18=> c0_n0_w18, 
            w19=> c0_n0_w19, 
            w20=> c0_n0_w20, 
            w21=> c0_n0_w21, 
            w22=> c0_n0_w22, 
            w23=> c0_n0_w23, 
            w24=> c0_n0_w24, 
            w25=> c0_n0_w25, 
            w26=> c0_n0_w26, 
            w27=> c0_n0_w27, 
            w28=> c0_n0_w28, 
            w29=> c0_n0_w29, 
            w30=> c0_n0_w30, 
            w31=> c0_n0_w31, 
            w32=> c0_n0_w32, 
            w33=> c0_n0_w33, 
            w34=> c0_n0_w34, 
            w35=> c0_n0_w35, 
            w36=> c0_n0_w36, 
            w37=> c0_n0_w37, 
            w38=> c0_n0_w38, 
            w39=> c0_n0_w39, 
            w40=> c0_n0_w40, 
            w41=> c0_n0_w41, 
            w42=> c0_n0_w42, 
            w43=> c0_n0_w43, 
            w44=> c0_n0_w44, 
            w45=> c0_n0_w45, 
            w46=> c0_n0_w46, 
            w47=> c0_n0_w47, 
            w48=> c0_n0_w48, 
            w49=> c0_n0_w49, 
            w50=> c0_n0_w50, 
            w51=> c0_n0_w51, 
            w52=> c0_n0_w52, 
            w53=> c0_n0_w53, 
            w54=> c0_n0_w54, 
            w55=> c0_n0_w55, 
            w56=> c0_n0_w56, 
            w57=> c0_n0_w57, 
            w58=> c0_n0_w58, 
            w59=> c0_n0_w59, 
            w60=> c0_n0_w60, 
            w61=> c0_n0_w61, 
            w62=> c0_n0_w62, 
            w63=> c0_n0_w63, 
            w64=> c0_n0_w64, 
            w65=> c0_n0_w65, 
            w66=> c0_n0_w66, 
            w67=> c0_n0_w67, 
            w68=> c0_n0_w68, 
            w69=> c0_n0_w69, 
            w70=> c0_n0_w70, 
            w71=> c0_n0_w71, 
            w72=> c0_n0_w72, 
            w73=> c0_n0_w73, 
            w74=> c0_n0_w74, 
            w75=> c0_n0_w75, 
            w76=> c0_n0_w76, 
            w77=> c0_n0_w77, 
            w78=> c0_n0_w78, 
            w79=> c0_n0_w79, 
            w80=> c0_n0_w80, 
            w81=> c0_n0_w81, 
            w82=> c0_n0_w82, 
            w83=> c0_n0_w83, 
            w84=> c0_n0_w84, 
            w85=> c0_n0_w85, 
            w86=> c0_n0_w86, 
            w87=> c0_n0_w87, 
            w88=> c0_n0_w88, 
            w89=> c0_n0_w89, 
            w90=> c0_n0_w90, 
            w91=> c0_n0_w91, 
            w92=> c0_n0_w92, 
            w93=> c0_n0_w93, 
            w94=> c0_n0_w94, 
            w95=> c0_n0_w95, 
            w96=> c0_n0_w96, 
            w97=> c0_n0_w97, 
            w98=> c0_n0_w98, 
            w99=> c0_n0_w99, 
            w100=> c0_n0_w100, 
            w101=> c0_n0_w101, 
            w102=> c0_n0_w102, 
            w103=> c0_n0_w103, 
            w104=> c0_n0_w104, 
            w105=> c0_n0_w105, 
            w106=> c0_n0_w106, 
            w107=> c0_n0_w107, 
            w108=> c0_n0_w108, 
            w109=> c0_n0_w109, 
            w110=> c0_n0_w110, 
            w111=> c0_n0_w111, 
            w112=> c0_n0_w112, 
            w113=> c0_n0_w113, 
            w114=> c0_n0_w114, 
            w115=> c0_n0_w115, 
            w116=> c0_n0_w116, 
            w117=> c0_n0_w117, 
            w118=> c0_n0_w118, 
            w119=> c0_n0_w119, 
            w120=> c0_n0_w120, 
            w121=> c0_n0_w121, 
            w122=> c0_n0_w122, 
            w123=> c0_n0_w123, 
            w124=> c0_n0_w124, 
            w125=> c0_n0_w125, 
            w126=> c0_n0_w126, 
            w127=> c0_n0_w127, 
            w128=> c0_n0_w128, 
            w129=> c0_n0_w129, 
            w130=> c0_n0_w130, 
            w131=> c0_n0_w131, 
            w132=> c0_n0_w132, 
            w133=> c0_n0_w133, 
            w134=> c0_n0_w134, 
            w135=> c0_n0_w135, 
            w136=> c0_n0_w136, 
            w137=> c0_n0_w137, 
            w138=> c0_n0_w138, 
            w139=> c0_n0_w139, 
            w140=> c0_n0_w140, 
            w141=> c0_n0_w141, 
            w142=> c0_n0_w142, 
            w143=> c0_n0_w143, 
            w144=> c0_n0_w144, 
            w145=> c0_n0_w145, 
            w146=> c0_n0_w146, 
            w147=> c0_n0_w147, 
            w148=> c0_n0_w148, 
            w149=> c0_n0_w149, 
            w150=> c0_n0_w150, 
            w151=> c0_n0_w151, 
            w152=> c0_n0_w152, 
            w153=> c0_n0_w153, 
            w154=> c0_n0_w154, 
            w155=> c0_n0_w155, 
            w156=> c0_n0_w156, 
            w157=> c0_n0_w157, 
            w158=> c0_n0_w158, 
            w159=> c0_n0_w159, 
            w160=> c0_n0_w160, 
            w161=> c0_n0_w161, 
            w162=> c0_n0_w162, 
            w163=> c0_n0_w163, 
            w164=> c0_n0_w164, 
            w165=> c0_n0_w165, 
            w166=> c0_n0_w166, 
            w167=> c0_n0_w167, 
            w168=> c0_n0_w168, 
            w169=> c0_n0_w169, 
            w170=> c0_n0_w170, 
            w171=> c0_n0_w171, 
            w172=> c0_n0_w172, 
            w173=> c0_n0_w173, 
            w174=> c0_n0_w174, 
            w175=> c0_n0_w175, 
            w176=> c0_n0_w176, 
            w177=> c0_n0_w177, 
            w178=> c0_n0_w178, 
            w179=> c0_n0_w179, 
            w180=> c0_n0_w180, 
            w181=> c0_n0_w181, 
            w182=> c0_n0_w182, 
            w183=> c0_n0_w183, 
            w184=> c0_n0_w184, 
            w185=> c0_n0_w185, 
            w186=> c0_n0_w186, 
            w187=> c0_n0_w187, 
            w188=> c0_n0_w188, 
            w189=> c0_n0_w189, 
            w190=> c0_n0_w190, 
            w191=> c0_n0_w191, 
            w192=> c0_n0_w192, 
            w193=> c0_n0_w193, 
            w194=> c0_n0_w194, 
            w195=> c0_n0_w195, 
            w196=> c0_n0_w196, 
            w197=> c0_n0_w197, 
            w198=> c0_n0_w198, 
            w199=> c0_n0_w199, 
            w200=> c0_n0_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n1_w1, 
            w2=> c0_n1_w2, 
            w3=> c0_n1_w3, 
            w4=> c0_n1_w4, 
            w5=> c0_n1_w5, 
            w6=> c0_n1_w6, 
            w7=> c0_n1_w7, 
            w8=> c0_n1_w8, 
            w9=> c0_n1_w9, 
            w10=> c0_n1_w10, 
            w11=> c0_n1_w11, 
            w12=> c0_n1_w12, 
            w13=> c0_n1_w13, 
            w14=> c0_n1_w14, 
            w15=> c0_n1_w15, 
            w16=> c0_n1_w16, 
            w17=> c0_n1_w17, 
            w18=> c0_n1_w18, 
            w19=> c0_n1_w19, 
            w20=> c0_n1_w20, 
            w21=> c0_n1_w21, 
            w22=> c0_n1_w22, 
            w23=> c0_n1_w23, 
            w24=> c0_n1_w24, 
            w25=> c0_n1_w25, 
            w26=> c0_n1_w26, 
            w27=> c0_n1_w27, 
            w28=> c0_n1_w28, 
            w29=> c0_n1_w29, 
            w30=> c0_n1_w30, 
            w31=> c0_n1_w31, 
            w32=> c0_n1_w32, 
            w33=> c0_n1_w33, 
            w34=> c0_n1_w34, 
            w35=> c0_n1_w35, 
            w36=> c0_n1_w36, 
            w37=> c0_n1_w37, 
            w38=> c0_n1_w38, 
            w39=> c0_n1_w39, 
            w40=> c0_n1_w40, 
            w41=> c0_n1_w41, 
            w42=> c0_n1_w42, 
            w43=> c0_n1_w43, 
            w44=> c0_n1_w44, 
            w45=> c0_n1_w45, 
            w46=> c0_n1_w46, 
            w47=> c0_n1_w47, 
            w48=> c0_n1_w48, 
            w49=> c0_n1_w49, 
            w50=> c0_n1_w50, 
            w51=> c0_n1_w51, 
            w52=> c0_n1_w52, 
            w53=> c0_n1_w53, 
            w54=> c0_n1_w54, 
            w55=> c0_n1_w55, 
            w56=> c0_n1_w56, 
            w57=> c0_n1_w57, 
            w58=> c0_n1_w58, 
            w59=> c0_n1_w59, 
            w60=> c0_n1_w60, 
            w61=> c0_n1_w61, 
            w62=> c0_n1_w62, 
            w63=> c0_n1_w63, 
            w64=> c0_n1_w64, 
            w65=> c0_n1_w65, 
            w66=> c0_n1_w66, 
            w67=> c0_n1_w67, 
            w68=> c0_n1_w68, 
            w69=> c0_n1_w69, 
            w70=> c0_n1_w70, 
            w71=> c0_n1_w71, 
            w72=> c0_n1_w72, 
            w73=> c0_n1_w73, 
            w74=> c0_n1_w74, 
            w75=> c0_n1_w75, 
            w76=> c0_n1_w76, 
            w77=> c0_n1_w77, 
            w78=> c0_n1_w78, 
            w79=> c0_n1_w79, 
            w80=> c0_n1_w80, 
            w81=> c0_n1_w81, 
            w82=> c0_n1_w82, 
            w83=> c0_n1_w83, 
            w84=> c0_n1_w84, 
            w85=> c0_n1_w85, 
            w86=> c0_n1_w86, 
            w87=> c0_n1_w87, 
            w88=> c0_n1_w88, 
            w89=> c0_n1_w89, 
            w90=> c0_n1_w90, 
            w91=> c0_n1_w91, 
            w92=> c0_n1_w92, 
            w93=> c0_n1_w93, 
            w94=> c0_n1_w94, 
            w95=> c0_n1_w95, 
            w96=> c0_n1_w96, 
            w97=> c0_n1_w97, 
            w98=> c0_n1_w98, 
            w99=> c0_n1_w99, 
            w100=> c0_n1_w100, 
            w101=> c0_n1_w101, 
            w102=> c0_n1_w102, 
            w103=> c0_n1_w103, 
            w104=> c0_n1_w104, 
            w105=> c0_n1_w105, 
            w106=> c0_n1_w106, 
            w107=> c0_n1_w107, 
            w108=> c0_n1_w108, 
            w109=> c0_n1_w109, 
            w110=> c0_n1_w110, 
            w111=> c0_n1_w111, 
            w112=> c0_n1_w112, 
            w113=> c0_n1_w113, 
            w114=> c0_n1_w114, 
            w115=> c0_n1_w115, 
            w116=> c0_n1_w116, 
            w117=> c0_n1_w117, 
            w118=> c0_n1_w118, 
            w119=> c0_n1_w119, 
            w120=> c0_n1_w120, 
            w121=> c0_n1_w121, 
            w122=> c0_n1_w122, 
            w123=> c0_n1_w123, 
            w124=> c0_n1_w124, 
            w125=> c0_n1_w125, 
            w126=> c0_n1_w126, 
            w127=> c0_n1_w127, 
            w128=> c0_n1_w128, 
            w129=> c0_n1_w129, 
            w130=> c0_n1_w130, 
            w131=> c0_n1_w131, 
            w132=> c0_n1_w132, 
            w133=> c0_n1_w133, 
            w134=> c0_n1_w134, 
            w135=> c0_n1_w135, 
            w136=> c0_n1_w136, 
            w137=> c0_n1_w137, 
            w138=> c0_n1_w138, 
            w139=> c0_n1_w139, 
            w140=> c0_n1_w140, 
            w141=> c0_n1_w141, 
            w142=> c0_n1_w142, 
            w143=> c0_n1_w143, 
            w144=> c0_n1_w144, 
            w145=> c0_n1_w145, 
            w146=> c0_n1_w146, 
            w147=> c0_n1_w147, 
            w148=> c0_n1_w148, 
            w149=> c0_n1_w149, 
            w150=> c0_n1_w150, 
            w151=> c0_n1_w151, 
            w152=> c0_n1_w152, 
            w153=> c0_n1_w153, 
            w154=> c0_n1_w154, 
            w155=> c0_n1_w155, 
            w156=> c0_n1_w156, 
            w157=> c0_n1_w157, 
            w158=> c0_n1_w158, 
            w159=> c0_n1_w159, 
            w160=> c0_n1_w160, 
            w161=> c0_n1_w161, 
            w162=> c0_n1_w162, 
            w163=> c0_n1_w163, 
            w164=> c0_n1_w164, 
            w165=> c0_n1_w165, 
            w166=> c0_n1_w166, 
            w167=> c0_n1_w167, 
            w168=> c0_n1_w168, 
            w169=> c0_n1_w169, 
            w170=> c0_n1_w170, 
            w171=> c0_n1_w171, 
            w172=> c0_n1_w172, 
            w173=> c0_n1_w173, 
            w174=> c0_n1_w174, 
            w175=> c0_n1_w175, 
            w176=> c0_n1_w176, 
            w177=> c0_n1_w177, 
            w178=> c0_n1_w178, 
            w179=> c0_n1_w179, 
            w180=> c0_n1_w180, 
            w181=> c0_n1_w181, 
            w182=> c0_n1_w182, 
            w183=> c0_n1_w183, 
            w184=> c0_n1_w184, 
            w185=> c0_n1_w185, 
            w186=> c0_n1_w186, 
            w187=> c0_n1_w187, 
            w188=> c0_n1_w188, 
            w189=> c0_n1_w189, 
            w190=> c0_n1_w190, 
            w191=> c0_n1_w191, 
            w192=> c0_n1_w192, 
            w193=> c0_n1_w193, 
            w194=> c0_n1_w194, 
            w195=> c0_n1_w195, 
            w196=> c0_n1_w196, 
            w197=> c0_n1_w197, 
            w198=> c0_n1_w198, 
            w199=> c0_n1_w199, 
            w200=> c0_n1_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n2_w1, 
            w2=> c0_n2_w2, 
            w3=> c0_n2_w3, 
            w4=> c0_n2_w4, 
            w5=> c0_n2_w5, 
            w6=> c0_n2_w6, 
            w7=> c0_n2_w7, 
            w8=> c0_n2_w8, 
            w9=> c0_n2_w9, 
            w10=> c0_n2_w10, 
            w11=> c0_n2_w11, 
            w12=> c0_n2_w12, 
            w13=> c0_n2_w13, 
            w14=> c0_n2_w14, 
            w15=> c0_n2_w15, 
            w16=> c0_n2_w16, 
            w17=> c0_n2_w17, 
            w18=> c0_n2_w18, 
            w19=> c0_n2_w19, 
            w20=> c0_n2_w20, 
            w21=> c0_n2_w21, 
            w22=> c0_n2_w22, 
            w23=> c0_n2_w23, 
            w24=> c0_n2_w24, 
            w25=> c0_n2_w25, 
            w26=> c0_n2_w26, 
            w27=> c0_n2_w27, 
            w28=> c0_n2_w28, 
            w29=> c0_n2_w29, 
            w30=> c0_n2_w30, 
            w31=> c0_n2_w31, 
            w32=> c0_n2_w32, 
            w33=> c0_n2_w33, 
            w34=> c0_n2_w34, 
            w35=> c0_n2_w35, 
            w36=> c0_n2_w36, 
            w37=> c0_n2_w37, 
            w38=> c0_n2_w38, 
            w39=> c0_n2_w39, 
            w40=> c0_n2_w40, 
            w41=> c0_n2_w41, 
            w42=> c0_n2_w42, 
            w43=> c0_n2_w43, 
            w44=> c0_n2_w44, 
            w45=> c0_n2_w45, 
            w46=> c0_n2_w46, 
            w47=> c0_n2_w47, 
            w48=> c0_n2_w48, 
            w49=> c0_n2_w49, 
            w50=> c0_n2_w50, 
            w51=> c0_n2_w51, 
            w52=> c0_n2_w52, 
            w53=> c0_n2_w53, 
            w54=> c0_n2_w54, 
            w55=> c0_n2_w55, 
            w56=> c0_n2_w56, 
            w57=> c0_n2_w57, 
            w58=> c0_n2_w58, 
            w59=> c0_n2_w59, 
            w60=> c0_n2_w60, 
            w61=> c0_n2_w61, 
            w62=> c0_n2_w62, 
            w63=> c0_n2_w63, 
            w64=> c0_n2_w64, 
            w65=> c0_n2_w65, 
            w66=> c0_n2_w66, 
            w67=> c0_n2_w67, 
            w68=> c0_n2_w68, 
            w69=> c0_n2_w69, 
            w70=> c0_n2_w70, 
            w71=> c0_n2_w71, 
            w72=> c0_n2_w72, 
            w73=> c0_n2_w73, 
            w74=> c0_n2_w74, 
            w75=> c0_n2_w75, 
            w76=> c0_n2_w76, 
            w77=> c0_n2_w77, 
            w78=> c0_n2_w78, 
            w79=> c0_n2_w79, 
            w80=> c0_n2_w80, 
            w81=> c0_n2_w81, 
            w82=> c0_n2_w82, 
            w83=> c0_n2_w83, 
            w84=> c0_n2_w84, 
            w85=> c0_n2_w85, 
            w86=> c0_n2_w86, 
            w87=> c0_n2_w87, 
            w88=> c0_n2_w88, 
            w89=> c0_n2_w89, 
            w90=> c0_n2_w90, 
            w91=> c0_n2_w91, 
            w92=> c0_n2_w92, 
            w93=> c0_n2_w93, 
            w94=> c0_n2_w94, 
            w95=> c0_n2_w95, 
            w96=> c0_n2_w96, 
            w97=> c0_n2_w97, 
            w98=> c0_n2_w98, 
            w99=> c0_n2_w99, 
            w100=> c0_n2_w100, 
            w101=> c0_n2_w101, 
            w102=> c0_n2_w102, 
            w103=> c0_n2_w103, 
            w104=> c0_n2_w104, 
            w105=> c0_n2_w105, 
            w106=> c0_n2_w106, 
            w107=> c0_n2_w107, 
            w108=> c0_n2_w108, 
            w109=> c0_n2_w109, 
            w110=> c0_n2_w110, 
            w111=> c0_n2_w111, 
            w112=> c0_n2_w112, 
            w113=> c0_n2_w113, 
            w114=> c0_n2_w114, 
            w115=> c0_n2_w115, 
            w116=> c0_n2_w116, 
            w117=> c0_n2_w117, 
            w118=> c0_n2_w118, 
            w119=> c0_n2_w119, 
            w120=> c0_n2_w120, 
            w121=> c0_n2_w121, 
            w122=> c0_n2_w122, 
            w123=> c0_n2_w123, 
            w124=> c0_n2_w124, 
            w125=> c0_n2_w125, 
            w126=> c0_n2_w126, 
            w127=> c0_n2_w127, 
            w128=> c0_n2_w128, 
            w129=> c0_n2_w129, 
            w130=> c0_n2_w130, 
            w131=> c0_n2_w131, 
            w132=> c0_n2_w132, 
            w133=> c0_n2_w133, 
            w134=> c0_n2_w134, 
            w135=> c0_n2_w135, 
            w136=> c0_n2_w136, 
            w137=> c0_n2_w137, 
            w138=> c0_n2_w138, 
            w139=> c0_n2_w139, 
            w140=> c0_n2_w140, 
            w141=> c0_n2_w141, 
            w142=> c0_n2_w142, 
            w143=> c0_n2_w143, 
            w144=> c0_n2_w144, 
            w145=> c0_n2_w145, 
            w146=> c0_n2_w146, 
            w147=> c0_n2_w147, 
            w148=> c0_n2_w148, 
            w149=> c0_n2_w149, 
            w150=> c0_n2_w150, 
            w151=> c0_n2_w151, 
            w152=> c0_n2_w152, 
            w153=> c0_n2_w153, 
            w154=> c0_n2_w154, 
            w155=> c0_n2_w155, 
            w156=> c0_n2_w156, 
            w157=> c0_n2_w157, 
            w158=> c0_n2_w158, 
            w159=> c0_n2_w159, 
            w160=> c0_n2_w160, 
            w161=> c0_n2_w161, 
            w162=> c0_n2_w162, 
            w163=> c0_n2_w163, 
            w164=> c0_n2_w164, 
            w165=> c0_n2_w165, 
            w166=> c0_n2_w166, 
            w167=> c0_n2_w167, 
            w168=> c0_n2_w168, 
            w169=> c0_n2_w169, 
            w170=> c0_n2_w170, 
            w171=> c0_n2_w171, 
            w172=> c0_n2_w172, 
            w173=> c0_n2_w173, 
            w174=> c0_n2_w174, 
            w175=> c0_n2_w175, 
            w176=> c0_n2_w176, 
            w177=> c0_n2_w177, 
            w178=> c0_n2_w178, 
            w179=> c0_n2_w179, 
            w180=> c0_n2_w180, 
            w181=> c0_n2_w181, 
            w182=> c0_n2_w182, 
            w183=> c0_n2_w183, 
            w184=> c0_n2_w184, 
            w185=> c0_n2_w185, 
            w186=> c0_n2_w186, 
            w187=> c0_n2_w187, 
            w188=> c0_n2_w188, 
            w189=> c0_n2_w189, 
            w190=> c0_n2_w190, 
            w191=> c0_n2_w191, 
            w192=> c0_n2_w192, 
            w193=> c0_n2_w193, 
            w194=> c0_n2_w194, 
            w195=> c0_n2_w195, 
            w196=> c0_n2_w196, 
            w197=> c0_n2_w197, 
            w198=> c0_n2_w198, 
            w199=> c0_n2_w199, 
            w200=> c0_n2_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n3_w1, 
            w2=> c0_n3_w2, 
            w3=> c0_n3_w3, 
            w4=> c0_n3_w4, 
            w5=> c0_n3_w5, 
            w6=> c0_n3_w6, 
            w7=> c0_n3_w7, 
            w8=> c0_n3_w8, 
            w9=> c0_n3_w9, 
            w10=> c0_n3_w10, 
            w11=> c0_n3_w11, 
            w12=> c0_n3_w12, 
            w13=> c0_n3_w13, 
            w14=> c0_n3_w14, 
            w15=> c0_n3_w15, 
            w16=> c0_n3_w16, 
            w17=> c0_n3_w17, 
            w18=> c0_n3_w18, 
            w19=> c0_n3_w19, 
            w20=> c0_n3_w20, 
            w21=> c0_n3_w21, 
            w22=> c0_n3_w22, 
            w23=> c0_n3_w23, 
            w24=> c0_n3_w24, 
            w25=> c0_n3_w25, 
            w26=> c0_n3_w26, 
            w27=> c0_n3_w27, 
            w28=> c0_n3_w28, 
            w29=> c0_n3_w29, 
            w30=> c0_n3_w30, 
            w31=> c0_n3_w31, 
            w32=> c0_n3_w32, 
            w33=> c0_n3_w33, 
            w34=> c0_n3_w34, 
            w35=> c0_n3_w35, 
            w36=> c0_n3_w36, 
            w37=> c0_n3_w37, 
            w38=> c0_n3_w38, 
            w39=> c0_n3_w39, 
            w40=> c0_n3_w40, 
            w41=> c0_n3_w41, 
            w42=> c0_n3_w42, 
            w43=> c0_n3_w43, 
            w44=> c0_n3_w44, 
            w45=> c0_n3_w45, 
            w46=> c0_n3_w46, 
            w47=> c0_n3_w47, 
            w48=> c0_n3_w48, 
            w49=> c0_n3_w49, 
            w50=> c0_n3_w50, 
            w51=> c0_n3_w51, 
            w52=> c0_n3_w52, 
            w53=> c0_n3_w53, 
            w54=> c0_n3_w54, 
            w55=> c0_n3_w55, 
            w56=> c0_n3_w56, 
            w57=> c0_n3_w57, 
            w58=> c0_n3_w58, 
            w59=> c0_n3_w59, 
            w60=> c0_n3_w60, 
            w61=> c0_n3_w61, 
            w62=> c0_n3_w62, 
            w63=> c0_n3_w63, 
            w64=> c0_n3_w64, 
            w65=> c0_n3_w65, 
            w66=> c0_n3_w66, 
            w67=> c0_n3_w67, 
            w68=> c0_n3_w68, 
            w69=> c0_n3_w69, 
            w70=> c0_n3_w70, 
            w71=> c0_n3_w71, 
            w72=> c0_n3_w72, 
            w73=> c0_n3_w73, 
            w74=> c0_n3_w74, 
            w75=> c0_n3_w75, 
            w76=> c0_n3_w76, 
            w77=> c0_n3_w77, 
            w78=> c0_n3_w78, 
            w79=> c0_n3_w79, 
            w80=> c0_n3_w80, 
            w81=> c0_n3_w81, 
            w82=> c0_n3_w82, 
            w83=> c0_n3_w83, 
            w84=> c0_n3_w84, 
            w85=> c0_n3_w85, 
            w86=> c0_n3_w86, 
            w87=> c0_n3_w87, 
            w88=> c0_n3_w88, 
            w89=> c0_n3_w89, 
            w90=> c0_n3_w90, 
            w91=> c0_n3_w91, 
            w92=> c0_n3_w92, 
            w93=> c0_n3_w93, 
            w94=> c0_n3_w94, 
            w95=> c0_n3_w95, 
            w96=> c0_n3_w96, 
            w97=> c0_n3_w97, 
            w98=> c0_n3_w98, 
            w99=> c0_n3_w99, 
            w100=> c0_n3_w100, 
            w101=> c0_n3_w101, 
            w102=> c0_n3_w102, 
            w103=> c0_n3_w103, 
            w104=> c0_n3_w104, 
            w105=> c0_n3_w105, 
            w106=> c0_n3_w106, 
            w107=> c0_n3_w107, 
            w108=> c0_n3_w108, 
            w109=> c0_n3_w109, 
            w110=> c0_n3_w110, 
            w111=> c0_n3_w111, 
            w112=> c0_n3_w112, 
            w113=> c0_n3_w113, 
            w114=> c0_n3_w114, 
            w115=> c0_n3_w115, 
            w116=> c0_n3_w116, 
            w117=> c0_n3_w117, 
            w118=> c0_n3_w118, 
            w119=> c0_n3_w119, 
            w120=> c0_n3_w120, 
            w121=> c0_n3_w121, 
            w122=> c0_n3_w122, 
            w123=> c0_n3_w123, 
            w124=> c0_n3_w124, 
            w125=> c0_n3_w125, 
            w126=> c0_n3_w126, 
            w127=> c0_n3_w127, 
            w128=> c0_n3_w128, 
            w129=> c0_n3_w129, 
            w130=> c0_n3_w130, 
            w131=> c0_n3_w131, 
            w132=> c0_n3_w132, 
            w133=> c0_n3_w133, 
            w134=> c0_n3_w134, 
            w135=> c0_n3_w135, 
            w136=> c0_n3_w136, 
            w137=> c0_n3_w137, 
            w138=> c0_n3_w138, 
            w139=> c0_n3_w139, 
            w140=> c0_n3_w140, 
            w141=> c0_n3_w141, 
            w142=> c0_n3_w142, 
            w143=> c0_n3_w143, 
            w144=> c0_n3_w144, 
            w145=> c0_n3_w145, 
            w146=> c0_n3_w146, 
            w147=> c0_n3_w147, 
            w148=> c0_n3_w148, 
            w149=> c0_n3_w149, 
            w150=> c0_n3_w150, 
            w151=> c0_n3_w151, 
            w152=> c0_n3_w152, 
            w153=> c0_n3_w153, 
            w154=> c0_n3_w154, 
            w155=> c0_n3_w155, 
            w156=> c0_n3_w156, 
            w157=> c0_n3_w157, 
            w158=> c0_n3_w158, 
            w159=> c0_n3_w159, 
            w160=> c0_n3_w160, 
            w161=> c0_n3_w161, 
            w162=> c0_n3_w162, 
            w163=> c0_n3_w163, 
            w164=> c0_n3_w164, 
            w165=> c0_n3_w165, 
            w166=> c0_n3_w166, 
            w167=> c0_n3_w167, 
            w168=> c0_n3_w168, 
            w169=> c0_n3_w169, 
            w170=> c0_n3_w170, 
            w171=> c0_n3_w171, 
            w172=> c0_n3_w172, 
            w173=> c0_n3_w173, 
            w174=> c0_n3_w174, 
            w175=> c0_n3_w175, 
            w176=> c0_n3_w176, 
            w177=> c0_n3_w177, 
            w178=> c0_n3_w178, 
            w179=> c0_n3_w179, 
            w180=> c0_n3_w180, 
            w181=> c0_n3_w181, 
            w182=> c0_n3_w182, 
            w183=> c0_n3_w183, 
            w184=> c0_n3_w184, 
            w185=> c0_n3_w185, 
            w186=> c0_n3_w186, 
            w187=> c0_n3_w187, 
            w188=> c0_n3_w188, 
            w189=> c0_n3_w189, 
            w190=> c0_n3_w190, 
            w191=> c0_n3_w191, 
            w192=> c0_n3_w192, 
            w193=> c0_n3_w193, 
            w194=> c0_n3_w194, 
            w195=> c0_n3_w195, 
            w196=> c0_n3_w196, 
            w197=> c0_n3_w197, 
            w198=> c0_n3_w198, 
            w199=> c0_n3_w199, 
            w200=> c0_n3_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n4_w1, 
            w2=> c0_n4_w2, 
            w3=> c0_n4_w3, 
            w4=> c0_n4_w4, 
            w5=> c0_n4_w5, 
            w6=> c0_n4_w6, 
            w7=> c0_n4_w7, 
            w8=> c0_n4_w8, 
            w9=> c0_n4_w9, 
            w10=> c0_n4_w10, 
            w11=> c0_n4_w11, 
            w12=> c0_n4_w12, 
            w13=> c0_n4_w13, 
            w14=> c0_n4_w14, 
            w15=> c0_n4_w15, 
            w16=> c0_n4_w16, 
            w17=> c0_n4_w17, 
            w18=> c0_n4_w18, 
            w19=> c0_n4_w19, 
            w20=> c0_n4_w20, 
            w21=> c0_n4_w21, 
            w22=> c0_n4_w22, 
            w23=> c0_n4_w23, 
            w24=> c0_n4_w24, 
            w25=> c0_n4_w25, 
            w26=> c0_n4_w26, 
            w27=> c0_n4_w27, 
            w28=> c0_n4_w28, 
            w29=> c0_n4_w29, 
            w30=> c0_n4_w30, 
            w31=> c0_n4_w31, 
            w32=> c0_n4_w32, 
            w33=> c0_n4_w33, 
            w34=> c0_n4_w34, 
            w35=> c0_n4_w35, 
            w36=> c0_n4_w36, 
            w37=> c0_n4_w37, 
            w38=> c0_n4_w38, 
            w39=> c0_n4_w39, 
            w40=> c0_n4_w40, 
            w41=> c0_n4_w41, 
            w42=> c0_n4_w42, 
            w43=> c0_n4_w43, 
            w44=> c0_n4_w44, 
            w45=> c0_n4_w45, 
            w46=> c0_n4_w46, 
            w47=> c0_n4_w47, 
            w48=> c0_n4_w48, 
            w49=> c0_n4_w49, 
            w50=> c0_n4_w50, 
            w51=> c0_n4_w51, 
            w52=> c0_n4_w52, 
            w53=> c0_n4_w53, 
            w54=> c0_n4_w54, 
            w55=> c0_n4_w55, 
            w56=> c0_n4_w56, 
            w57=> c0_n4_w57, 
            w58=> c0_n4_w58, 
            w59=> c0_n4_w59, 
            w60=> c0_n4_w60, 
            w61=> c0_n4_w61, 
            w62=> c0_n4_w62, 
            w63=> c0_n4_w63, 
            w64=> c0_n4_w64, 
            w65=> c0_n4_w65, 
            w66=> c0_n4_w66, 
            w67=> c0_n4_w67, 
            w68=> c0_n4_w68, 
            w69=> c0_n4_w69, 
            w70=> c0_n4_w70, 
            w71=> c0_n4_w71, 
            w72=> c0_n4_w72, 
            w73=> c0_n4_w73, 
            w74=> c0_n4_w74, 
            w75=> c0_n4_w75, 
            w76=> c0_n4_w76, 
            w77=> c0_n4_w77, 
            w78=> c0_n4_w78, 
            w79=> c0_n4_w79, 
            w80=> c0_n4_w80, 
            w81=> c0_n4_w81, 
            w82=> c0_n4_w82, 
            w83=> c0_n4_w83, 
            w84=> c0_n4_w84, 
            w85=> c0_n4_w85, 
            w86=> c0_n4_w86, 
            w87=> c0_n4_w87, 
            w88=> c0_n4_w88, 
            w89=> c0_n4_w89, 
            w90=> c0_n4_w90, 
            w91=> c0_n4_w91, 
            w92=> c0_n4_w92, 
            w93=> c0_n4_w93, 
            w94=> c0_n4_w94, 
            w95=> c0_n4_w95, 
            w96=> c0_n4_w96, 
            w97=> c0_n4_w97, 
            w98=> c0_n4_w98, 
            w99=> c0_n4_w99, 
            w100=> c0_n4_w100, 
            w101=> c0_n4_w101, 
            w102=> c0_n4_w102, 
            w103=> c0_n4_w103, 
            w104=> c0_n4_w104, 
            w105=> c0_n4_w105, 
            w106=> c0_n4_w106, 
            w107=> c0_n4_w107, 
            w108=> c0_n4_w108, 
            w109=> c0_n4_w109, 
            w110=> c0_n4_w110, 
            w111=> c0_n4_w111, 
            w112=> c0_n4_w112, 
            w113=> c0_n4_w113, 
            w114=> c0_n4_w114, 
            w115=> c0_n4_w115, 
            w116=> c0_n4_w116, 
            w117=> c0_n4_w117, 
            w118=> c0_n4_w118, 
            w119=> c0_n4_w119, 
            w120=> c0_n4_w120, 
            w121=> c0_n4_w121, 
            w122=> c0_n4_w122, 
            w123=> c0_n4_w123, 
            w124=> c0_n4_w124, 
            w125=> c0_n4_w125, 
            w126=> c0_n4_w126, 
            w127=> c0_n4_w127, 
            w128=> c0_n4_w128, 
            w129=> c0_n4_w129, 
            w130=> c0_n4_w130, 
            w131=> c0_n4_w131, 
            w132=> c0_n4_w132, 
            w133=> c0_n4_w133, 
            w134=> c0_n4_w134, 
            w135=> c0_n4_w135, 
            w136=> c0_n4_w136, 
            w137=> c0_n4_w137, 
            w138=> c0_n4_w138, 
            w139=> c0_n4_w139, 
            w140=> c0_n4_w140, 
            w141=> c0_n4_w141, 
            w142=> c0_n4_w142, 
            w143=> c0_n4_w143, 
            w144=> c0_n4_w144, 
            w145=> c0_n4_w145, 
            w146=> c0_n4_w146, 
            w147=> c0_n4_w147, 
            w148=> c0_n4_w148, 
            w149=> c0_n4_w149, 
            w150=> c0_n4_w150, 
            w151=> c0_n4_w151, 
            w152=> c0_n4_w152, 
            w153=> c0_n4_w153, 
            w154=> c0_n4_w154, 
            w155=> c0_n4_w155, 
            w156=> c0_n4_w156, 
            w157=> c0_n4_w157, 
            w158=> c0_n4_w158, 
            w159=> c0_n4_w159, 
            w160=> c0_n4_w160, 
            w161=> c0_n4_w161, 
            w162=> c0_n4_w162, 
            w163=> c0_n4_w163, 
            w164=> c0_n4_w164, 
            w165=> c0_n4_w165, 
            w166=> c0_n4_w166, 
            w167=> c0_n4_w167, 
            w168=> c0_n4_w168, 
            w169=> c0_n4_w169, 
            w170=> c0_n4_w170, 
            w171=> c0_n4_w171, 
            w172=> c0_n4_w172, 
            w173=> c0_n4_w173, 
            w174=> c0_n4_w174, 
            w175=> c0_n4_w175, 
            w176=> c0_n4_w176, 
            w177=> c0_n4_w177, 
            w178=> c0_n4_w178, 
            w179=> c0_n4_w179, 
            w180=> c0_n4_w180, 
            w181=> c0_n4_w181, 
            w182=> c0_n4_w182, 
            w183=> c0_n4_w183, 
            w184=> c0_n4_w184, 
            w185=> c0_n4_w185, 
            w186=> c0_n4_w186, 
            w187=> c0_n4_w187, 
            w188=> c0_n4_w188, 
            w189=> c0_n4_w189, 
            w190=> c0_n4_w190, 
            w191=> c0_n4_w191, 
            w192=> c0_n4_w192, 
            w193=> c0_n4_w193, 
            w194=> c0_n4_w194, 
            w195=> c0_n4_w195, 
            w196=> c0_n4_w196, 
            w197=> c0_n4_w197, 
            w198=> c0_n4_w198, 
            w199=> c0_n4_w199, 
            w200=> c0_n4_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n5_w1, 
            w2=> c0_n5_w2, 
            w3=> c0_n5_w3, 
            w4=> c0_n5_w4, 
            w5=> c0_n5_w5, 
            w6=> c0_n5_w6, 
            w7=> c0_n5_w7, 
            w8=> c0_n5_w8, 
            w9=> c0_n5_w9, 
            w10=> c0_n5_w10, 
            w11=> c0_n5_w11, 
            w12=> c0_n5_w12, 
            w13=> c0_n5_w13, 
            w14=> c0_n5_w14, 
            w15=> c0_n5_w15, 
            w16=> c0_n5_w16, 
            w17=> c0_n5_w17, 
            w18=> c0_n5_w18, 
            w19=> c0_n5_w19, 
            w20=> c0_n5_w20, 
            w21=> c0_n5_w21, 
            w22=> c0_n5_w22, 
            w23=> c0_n5_w23, 
            w24=> c0_n5_w24, 
            w25=> c0_n5_w25, 
            w26=> c0_n5_w26, 
            w27=> c0_n5_w27, 
            w28=> c0_n5_w28, 
            w29=> c0_n5_w29, 
            w30=> c0_n5_w30, 
            w31=> c0_n5_w31, 
            w32=> c0_n5_w32, 
            w33=> c0_n5_w33, 
            w34=> c0_n5_w34, 
            w35=> c0_n5_w35, 
            w36=> c0_n5_w36, 
            w37=> c0_n5_w37, 
            w38=> c0_n5_w38, 
            w39=> c0_n5_w39, 
            w40=> c0_n5_w40, 
            w41=> c0_n5_w41, 
            w42=> c0_n5_w42, 
            w43=> c0_n5_w43, 
            w44=> c0_n5_w44, 
            w45=> c0_n5_w45, 
            w46=> c0_n5_w46, 
            w47=> c0_n5_w47, 
            w48=> c0_n5_w48, 
            w49=> c0_n5_w49, 
            w50=> c0_n5_w50, 
            w51=> c0_n5_w51, 
            w52=> c0_n5_w52, 
            w53=> c0_n5_w53, 
            w54=> c0_n5_w54, 
            w55=> c0_n5_w55, 
            w56=> c0_n5_w56, 
            w57=> c0_n5_w57, 
            w58=> c0_n5_w58, 
            w59=> c0_n5_w59, 
            w60=> c0_n5_w60, 
            w61=> c0_n5_w61, 
            w62=> c0_n5_w62, 
            w63=> c0_n5_w63, 
            w64=> c0_n5_w64, 
            w65=> c0_n5_w65, 
            w66=> c0_n5_w66, 
            w67=> c0_n5_w67, 
            w68=> c0_n5_w68, 
            w69=> c0_n5_w69, 
            w70=> c0_n5_w70, 
            w71=> c0_n5_w71, 
            w72=> c0_n5_w72, 
            w73=> c0_n5_w73, 
            w74=> c0_n5_w74, 
            w75=> c0_n5_w75, 
            w76=> c0_n5_w76, 
            w77=> c0_n5_w77, 
            w78=> c0_n5_w78, 
            w79=> c0_n5_w79, 
            w80=> c0_n5_w80, 
            w81=> c0_n5_w81, 
            w82=> c0_n5_w82, 
            w83=> c0_n5_w83, 
            w84=> c0_n5_w84, 
            w85=> c0_n5_w85, 
            w86=> c0_n5_w86, 
            w87=> c0_n5_w87, 
            w88=> c0_n5_w88, 
            w89=> c0_n5_w89, 
            w90=> c0_n5_w90, 
            w91=> c0_n5_w91, 
            w92=> c0_n5_w92, 
            w93=> c0_n5_w93, 
            w94=> c0_n5_w94, 
            w95=> c0_n5_w95, 
            w96=> c0_n5_w96, 
            w97=> c0_n5_w97, 
            w98=> c0_n5_w98, 
            w99=> c0_n5_w99, 
            w100=> c0_n5_w100, 
            w101=> c0_n5_w101, 
            w102=> c0_n5_w102, 
            w103=> c0_n5_w103, 
            w104=> c0_n5_w104, 
            w105=> c0_n5_w105, 
            w106=> c0_n5_w106, 
            w107=> c0_n5_w107, 
            w108=> c0_n5_w108, 
            w109=> c0_n5_w109, 
            w110=> c0_n5_w110, 
            w111=> c0_n5_w111, 
            w112=> c0_n5_w112, 
            w113=> c0_n5_w113, 
            w114=> c0_n5_w114, 
            w115=> c0_n5_w115, 
            w116=> c0_n5_w116, 
            w117=> c0_n5_w117, 
            w118=> c0_n5_w118, 
            w119=> c0_n5_w119, 
            w120=> c0_n5_w120, 
            w121=> c0_n5_w121, 
            w122=> c0_n5_w122, 
            w123=> c0_n5_w123, 
            w124=> c0_n5_w124, 
            w125=> c0_n5_w125, 
            w126=> c0_n5_w126, 
            w127=> c0_n5_w127, 
            w128=> c0_n5_w128, 
            w129=> c0_n5_w129, 
            w130=> c0_n5_w130, 
            w131=> c0_n5_w131, 
            w132=> c0_n5_w132, 
            w133=> c0_n5_w133, 
            w134=> c0_n5_w134, 
            w135=> c0_n5_w135, 
            w136=> c0_n5_w136, 
            w137=> c0_n5_w137, 
            w138=> c0_n5_w138, 
            w139=> c0_n5_w139, 
            w140=> c0_n5_w140, 
            w141=> c0_n5_w141, 
            w142=> c0_n5_w142, 
            w143=> c0_n5_w143, 
            w144=> c0_n5_w144, 
            w145=> c0_n5_w145, 
            w146=> c0_n5_w146, 
            w147=> c0_n5_w147, 
            w148=> c0_n5_w148, 
            w149=> c0_n5_w149, 
            w150=> c0_n5_w150, 
            w151=> c0_n5_w151, 
            w152=> c0_n5_w152, 
            w153=> c0_n5_w153, 
            w154=> c0_n5_w154, 
            w155=> c0_n5_w155, 
            w156=> c0_n5_w156, 
            w157=> c0_n5_w157, 
            w158=> c0_n5_w158, 
            w159=> c0_n5_w159, 
            w160=> c0_n5_w160, 
            w161=> c0_n5_w161, 
            w162=> c0_n5_w162, 
            w163=> c0_n5_w163, 
            w164=> c0_n5_w164, 
            w165=> c0_n5_w165, 
            w166=> c0_n5_w166, 
            w167=> c0_n5_w167, 
            w168=> c0_n5_w168, 
            w169=> c0_n5_w169, 
            w170=> c0_n5_w170, 
            w171=> c0_n5_w171, 
            w172=> c0_n5_w172, 
            w173=> c0_n5_w173, 
            w174=> c0_n5_w174, 
            w175=> c0_n5_w175, 
            w176=> c0_n5_w176, 
            w177=> c0_n5_w177, 
            w178=> c0_n5_w178, 
            w179=> c0_n5_w179, 
            w180=> c0_n5_w180, 
            w181=> c0_n5_w181, 
            w182=> c0_n5_w182, 
            w183=> c0_n5_w183, 
            w184=> c0_n5_w184, 
            w185=> c0_n5_w185, 
            w186=> c0_n5_w186, 
            w187=> c0_n5_w187, 
            w188=> c0_n5_w188, 
            w189=> c0_n5_w189, 
            w190=> c0_n5_w190, 
            w191=> c0_n5_w191, 
            w192=> c0_n5_w192, 
            w193=> c0_n5_w193, 
            w194=> c0_n5_w194, 
            w195=> c0_n5_w195, 
            w196=> c0_n5_w196, 
            w197=> c0_n5_w197, 
            w198=> c0_n5_w198, 
            w199=> c0_n5_w199, 
            w200=> c0_n5_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n6_w1, 
            w2=> c0_n6_w2, 
            w3=> c0_n6_w3, 
            w4=> c0_n6_w4, 
            w5=> c0_n6_w5, 
            w6=> c0_n6_w6, 
            w7=> c0_n6_w7, 
            w8=> c0_n6_w8, 
            w9=> c0_n6_w9, 
            w10=> c0_n6_w10, 
            w11=> c0_n6_w11, 
            w12=> c0_n6_w12, 
            w13=> c0_n6_w13, 
            w14=> c0_n6_w14, 
            w15=> c0_n6_w15, 
            w16=> c0_n6_w16, 
            w17=> c0_n6_w17, 
            w18=> c0_n6_w18, 
            w19=> c0_n6_w19, 
            w20=> c0_n6_w20, 
            w21=> c0_n6_w21, 
            w22=> c0_n6_w22, 
            w23=> c0_n6_w23, 
            w24=> c0_n6_w24, 
            w25=> c0_n6_w25, 
            w26=> c0_n6_w26, 
            w27=> c0_n6_w27, 
            w28=> c0_n6_w28, 
            w29=> c0_n6_w29, 
            w30=> c0_n6_w30, 
            w31=> c0_n6_w31, 
            w32=> c0_n6_w32, 
            w33=> c0_n6_w33, 
            w34=> c0_n6_w34, 
            w35=> c0_n6_w35, 
            w36=> c0_n6_w36, 
            w37=> c0_n6_w37, 
            w38=> c0_n6_w38, 
            w39=> c0_n6_w39, 
            w40=> c0_n6_w40, 
            w41=> c0_n6_w41, 
            w42=> c0_n6_w42, 
            w43=> c0_n6_w43, 
            w44=> c0_n6_w44, 
            w45=> c0_n6_w45, 
            w46=> c0_n6_w46, 
            w47=> c0_n6_w47, 
            w48=> c0_n6_w48, 
            w49=> c0_n6_w49, 
            w50=> c0_n6_w50, 
            w51=> c0_n6_w51, 
            w52=> c0_n6_w52, 
            w53=> c0_n6_w53, 
            w54=> c0_n6_w54, 
            w55=> c0_n6_w55, 
            w56=> c0_n6_w56, 
            w57=> c0_n6_w57, 
            w58=> c0_n6_w58, 
            w59=> c0_n6_w59, 
            w60=> c0_n6_w60, 
            w61=> c0_n6_w61, 
            w62=> c0_n6_w62, 
            w63=> c0_n6_w63, 
            w64=> c0_n6_w64, 
            w65=> c0_n6_w65, 
            w66=> c0_n6_w66, 
            w67=> c0_n6_w67, 
            w68=> c0_n6_w68, 
            w69=> c0_n6_w69, 
            w70=> c0_n6_w70, 
            w71=> c0_n6_w71, 
            w72=> c0_n6_w72, 
            w73=> c0_n6_w73, 
            w74=> c0_n6_w74, 
            w75=> c0_n6_w75, 
            w76=> c0_n6_w76, 
            w77=> c0_n6_w77, 
            w78=> c0_n6_w78, 
            w79=> c0_n6_w79, 
            w80=> c0_n6_w80, 
            w81=> c0_n6_w81, 
            w82=> c0_n6_w82, 
            w83=> c0_n6_w83, 
            w84=> c0_n6_w84, 
            w85=> c0_n6_w85, 
            w86=> c0_n6_w86, 
            w87=> c0_n6_w87, 
            w88=> c0_n6_w88, 
            w89=> c0_n6_w89, 
            w90=> c0_n6_w90, 
            w91=> c0_n6_w91, 
            w92=> c0_n6_w92, 
            w93=> c0_n6_w93, 
            w94=> c0_n6_w94, 
            w95=> c0_n6_w95, 
            w96=> c0_n6_w96, 
            w97=> c0_n6_w97, 
            w98=> c0_n6_w98, 
            w99=> c0_n6_w99, 
            w100=> c0_n6_w100, 
            w101=> c0_n6_w101, 
            w102=> c0_n6_w102, 
            w103=> c0_n6_w103, 
            w104=> c0_n6_w104, 
            w105=> c0_n6_w105, 
            w106=> c0_n6_w106, 
            w107=> c0_n6_w107, 
            w108=> c0_n6_w108, 
            w109=> c0_n6_w109, 
            w110=> c0_n6_w110, 
            w111=> c0_n6_w111, 
            w112=> c0_n6_w112, 
            w113=> c0_n6_w113, 
            w114=> c0_n6_w114, 
            w115=> c0_n6_w115, 
            w116=> c0_n6_w116, 
            w117=> c0_n6_w117, 
            w118=> c0_n6_w118, 
            w119=> c0_n6_w119, 
            w120=> c0_n6_w120, 
            w121=> c0_n6_w121, 
            w122=> c0_n6_w122, 
            w123=> c0_n6_w123, 
            w124=> c0_n6_w124, 
            w125=> c0_n6_w125, 
            w126=> c0_n6_w126, 
            w127=> c0_n6_w127, 
            w128=> c0_n6_w128, 
            w129=> c0_n6_w129, 
            w130=> c0_n6_w130, 
            w131=> c0_n6_w131, 
            w132=> c0_n6_w132, 
            w133=> c0_n6_w133, 
            w134=> c0_n6_w134, 
            w135=> c0_n6_w135, 
            w136=> c0_n6_w136, 
            w137=> c0_n6_w137, 
            w138=> c0_n6_w138, 
            w139=> c0_n6_w139, 
            w140=> c0_n6_w140, 
            w141=> c0_n6_w141, 
            w142=> c0_n6_w142, 
            w143=> c0_n6_w143, 
            w144=> c0_n6_w144, 
            w145=> c0_n6_w145, 
            w146=> c0_n6_w146, 
            w147=> c0_n6_w147, 
            w148=> c0_n6_w148, 
            w149=> c0_n6_w149, 
            w150=> c0_n6_w150, 
            w151=> c0_n6_w151, 
            w152=> c0_n6_w152, 
            w153=> c0_n6_w153, 
            w154=> c0_n6_w154, 
            w155=> c0_n6_w155, 
            w156=> c0_n6_w156, 
            w157=> c0_n6_w157, 
            w158=> c0_n6_w158, 
            w159=> c0_n6_w159, 
            w160=> c0_n6_w160, 
            w161=> c0_n6_w161, 
            w162=> c0_n6_w162, 
            w163=> c0_n6_w163, 
            w164=> c0_n6_w164, 
            w165=> c0_n6_w165, 
            w166=> c0_n6_w166, 
            w167=> c0_n6_w167, 
            w168=> c0_n6_w168, 
            w169=> c0_n6_w169, 
            w170=> c0_n6_w170, 
            w171=> c0_n6_w171, 
            w172=> c0_n6_w172, 
            w173=> c0_n6_w173, 
            w174=> c0_n6_w174, 
            w175=> c0_n6_w175, 
            w176=> c0_n6_w176, 
            w177=> c0_n6_w177, 
            w178=> c0_n6_w178, 
            w179=> c0_n6_w179, 
            w180=> c0_n6_w180, 
            w181=> c0_n6_w181, 
            w182=> c0_n6_w182, 
            w183=> c0_n6_w183, 
            w184=> c0_n6_w184, 
            w185=> c0_n6_w185, 
            w186=> c0_n6_w186, 
            w187=> c0_n6_w187, 
            w188=> c0_n6_w188, 
            w189=> c0_n6_w189, 
            w190=> c0_n6_w190, 
            w191=> c0_n6_w191, 
            w192=> c0_n6_w192, 
            w193=> c0_n6_w193, 
            w194=> c0_n6_w194, 
            w195=> c0_n6_w195, 
            w196=> c0_n6_w196, 
            w197=> c0_n6_w197, 
            w198=> c0_n6_w198, 
            w199=> c0_n6_w199, 
            w200=> c0_n6_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n7_w1, 
            w2=> c0_n7_w2, 
            w3=> c0_n7_w3, 
            w4=> c0_n7_w4, 
            w5=> c0_n7_w5, 
            w6=> c0_n7_w6, 
            w7=> c0_n7_w7, 
            w8=> c0_n7_w8, 
            w9=> c0_n7_w9, 
            w10=> c0_n7_w10, 
            w11=> c0_n7_w11, 
            w12=> c0_n7_w12, 
            w13=> c0_n7_w13, 
            w14=> c0_n7_w14, 
            w15=> c0_n7_w15, 
            w16=> c0_n7_w16, 
            w17=> c0_n7_w17, 
            w18=> c0_n7_w18, 
            w19=> c0_n7_w19, 
            w20=> c0_n7_w20, 
            w21=> c0_n7_w21, 
            w22=> c0_n7_w22, 
            w23=> c0_n7_w23, 
            w24=> c0_n7_w24, 
            w25=> c0_n7_w25, 
            w26=> c0_n7_w26, 
            w27=> c0_n7_w27, 
            w28=> c0_n7_w28, 
            w29=> c0_n7_w29, 
            w30=> c0_n7_w30, 
            w31=> c0_n7_w31, 
            w32=> c0_n7_w32, 
            w33=> c0_n7_w33, 
            w34=> c0_n7_w34, 
            w35=> c0_n7_w35, 
            w36=> c0_n7_w36, 
            w37=> c0_n7_w37, 
            w38=> c0_n7_w38, 
            w39=> c0_n7_w39, 
            w40=> c0_n7_w40, 
            w41=> c0_n7_w41, 
            w42=> c0_n7_w42, 
            w43=> c0_n7_w43, 
            w44=> c0_n7_w44, 
            w45=> c0_n7_w45, 
            w46=> c0_n7_w46, 
            w47=> c0_n7_w47, 
            w48=> c0_n7_w48, 
            w49=> c0_n7_w49, 
            w50=> c0_n7_w50, 
            w51=> c0_n7_w51, 
            w52=> c0_n7_w52, 
            w53=> c0_n7_w53, 
            w54=> c0_n7_w54, 
            w55=> c0_n7_w55, 
            w56=> c0_n7_w56, 
            w57=> c0_n7_w57, 
            w58=> c0_n7_w58, 
            w59=> c0_n7_w59, 
            w60=> c0_n7_w60, 
            w61=> c0_n7_w61, 
            w62=> c0_n7_w62, 
            w63=> c0_n7_w63, 
            w64=> c0_n7_w64, 
            w65=> c0_n7_w65, 
            w66=> c0_n7_w66, 
            w67=> c0_n7_w67, 
            w68=> c0_n7_w68, 
            w69=> c0_n7_w69, 
            w70=> c0_n7_w70, 
            w71=> c0_n7_w71, 
            w72=> c0_n7_w72, 
            w73=> c0_n7_w73, 
            w74=> c0_n7_w74, 
            w75=> c0_n7_w75, 
            w76=> c0_n7_w76, 
            w77=> c0_n7_w77, 
            w78=> c0_n7_w78, 
            w79=> c0_n7_w79, 
            w80=> c0_n7_w80, 
            w81=> c0_n7_w81, 
            w82=> c0_n7_w82, 
            w83=> c0_n7_w83, 
            w84=> c0_n7_w84, 
            w85=> c0_n7_w85, 
            w86=> c0_n7_w86, 
            w87=> c0_n7_w87, 
            w88=> c0_n7_w88, 
            w89=> c0_n7_w89, 
            w90=> c0_n7_w90, 
            w91=> c0_n7_w91, 
            w92=> c0_n7_w92, 
            w93=> c0_n7_w93, 
            w94=> c0_n7_w94, 
            w95=> c0_n7_w95, 
            w96=> c0_n7_w96, 
            w97=> c0_n7_w97, 
            w98=> c0_n7_w98, 
            w99=> c0_n7_w99, 
            w100=> c0_n7_w100, 
            w101=> c0_n7_w101, 
            w102=> c0_n7_w102, 
            w103=> c0_n7_w103, 
            w104=> c0_n7_w104, 
            w105=> c0_n7_w105, 
            w106=> c0_n7_w106, 
            w107=> c0_n7_w107, 
            w108=> c0_n7_w108, 
            w109=> c0_n7_w109, 
            w110=> c0_n7_w110, 
            w111=> c0_n7_w111, 
            w112=> c0_n7_w112, 
            w113=> c0_n7_w113, 
            w114=> c0_n7_w114, 
            w115=> c0_n7_w115, 
            w116=> c0_n7_w116, 
            w117=> c0_n7_w117, 
            w118=> c0_n7_w118, 
            w119=> c0_n7_w119, 
            w120=> c0_n7_w120, 
            w121=> c0_n7_w121, 
            w122=> c0_n7_w122, 
            w123=> c0_n7_w123, 
            w124=> c0_n7_w124, 
            w125=> c0_n7_w125, 
            w126=> c0_n7_w126, 
            w127=> c0_n7_w127, 
            w128=> c0_n7_w128, 
            w129=> c0_n7_w129, 
            w130=> c0_n7_w130, 
            w131=> c0_n7_w131, 
            w132=> c0_n7_w132, 
            w133=> c0_n7_w133, 
            w134=> c0_n7_w134, 
            w135=> c0_n7_w135, 
            w136=> c0_n7_w136, 
            w137=> c0_n7_w137, 
            w138=> c0_n7_w138, 
            w139=> c0_n7_w139, 
            w140=> c0_n7_w140, 
            w141=> c0_n7_w141, 
            w142=> c0_n7_w142, 
            w143=> c0_n7_w143, 
            w144=> c0_n7_w144, 
            w145=> c0_n7_w145, 
            w146=> c0_n7_w146, 
            w147=> c0_n7_w147, 
            w148=> c0_n7_w148, 
            w149=> c0_n7_w149, 
            w150=> c0_n7_w150, 
            w151=> c0_n7_w151, 
            w152=> c0_n7_w152, 
            w153=> c0_n7_w153, 
            w154=> c0_n7_w154, 
            w155=> c0_n7_w155, 
            w156=> c0_n7_w156, 
            w157=> c0_n7_w157, 
            w158=> c0_n7_w158, 
            w159=> c0_n7_w159, 
            w160=> c0_n7_w160, 
            w161=> c0_n7_w161, 
            w162=> c0_n7_w162, 
            w163=> c0_n7_w163, 
            w164=> c0_n7_w164, 
            w165=> c0_n7_w165, 
            w166=> c0_n7_w166, 
            w167=> c0_n7_w167, 
            w168=> c0_n7_w168, 
            w169=> c0_n7_w169, 
            w170=> c0_n7_w170, 
            w171=> c0_n7_w171, 
            w172=> c0_n7_w172, 
            w173=> c0_n7_w173, 
            w174=> c0_n7_w174, 
            w175=> c0_n7_w175, 
            w176=> c0_n7_w176, 
            w177=> c0_n7_w177, 
            w178=> c0_n7_w178, 
            w179=> c0_n7_w179, 
            w180=> c0_n7_w180, 
            w181=> c0_n7_w181, 
            w182=> c0_n7_w182, 
            w183=> c0_n7_w183, 
            w184=> c0_n7_w184, 
            w185=> c0_n7_w185, 
            w186=> c0_n7_w186, 
            w187=> c0_n7_w187, 
            w188=> c0_n7_w188, 
            w189=> c0_n7_w189, 
            w190=> c0_n7_w190, 
            w191=> c0_n7_w191, 
            w192=> c0_n7_w192, 
            w193=> c0_n7_w193, 
            w194=> c0_n7_w194, 
            w195=> c0_n7_w195, 
            w196=> c0_n7_w196, 
            w197=> c0_n7_w197, 
            w198=> c0_n7_w198, 
            w199=> c0_n7_w199, 
            w200=> c0_n7_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n8_w1, 
            w2=> c0_n8_w2, 
            w3=> c0_n8_w3, 
            w4=> c0_n8_w4, 
            w5=> c0_n8_w5, 
            w6=> c0_n8_w6, 
            w7=> c0_n8_w7, 
            w8=> c0_n8_w8, 
            w9=> c0_n8_w9, 
            w10=> c0_n8_w10, 
            w11=> c0_n8_w11, 
            w12=> c0_n8_w12, 
            w13=> c0_n8_w13, 
            w14=> c0_n8_w14, 
            w15=> c0_n8_w15, 
            w16=> c0_n8_w16, 
            w17=> c0_n8_w17, 
            w18=> c0_n8_w18, 
            w19=> c0_n8_w19, 
            w20=> c0_n8_w20, 
            w21=> c0_n8_w21, 
            w22=> c0_n8_w22, 
            w23=> c0_n8_w23, 
            w24=> c0_n8_w24, 
            w25=> c0_n8_w25, 
            w26=> c0_n8_w26, 
            w27=> c0_n8_w27, 
            w28=> c0_n8_w28, 
            w29=> c0_n8_w29, 
            w30=> c0_n8_w30, 
            w31=> c0_n8_w31, 
            w32=> c0_n8_w32, 
            w33=> c0_n8_w33, 
            w34=> c0_n8_w34, 
            w35=> c0_n8_w35, 
            w36=> c0_n8_w36, 
            w37=> c0_n8_w37, 
            w38=> c0_n8_w38, 
            w39=> c0_n8_w39, 
            w40=> c0_n8_w40, 
            w41=> c0_n8_w41, 
            w42=> c0_n8_w42, 
            w43=> c0_n8_w43, 
            w44=> c0_n8_w44, 
            w45=> c0_n8_w45, 
            w46=> c0_n8_w46, 
            w47=> c0_n8_w47, 
            w48=> c0_n8_w48, 
            w49=> c0_n8_w49, 
            w50=> c0_n8_w50, 
            w51=> c0_n8_w51, 
            w52=> c0_n8_w52, 
            w53=> c0_n8_w53, 
            w54=> c0_n8_w54, 
            w55=> c0_n8_w55, 
            w56=> c0_n8_w56, 
            w57=> c0_n8_w57, 
            w58=> c0_n8_w58, 
            w59=> c0_n8_w59, 
            w60=> c0_n8_w60, 
            w61=> c0_n8_w61, 
            w62=> c0_n8_w62, 
            w63=> c0_n8_w63, 
            w64=> c0_n8_w64, 
            w65=> c0_n8_w65, 
            w66=> c0_n8_w66, 
            w67=> c0_n8_w67, 
            w68=> c0_n8_w68, 
            w69=> c0_n8_w69, 
            w70=> c0_n8_w70, 
            w71=> c0_n8_w71, 
            w72=> c0_n8_w72, 
            w73=> c0_n8_w73, 
            w74=> c0_n8_w74, 
            w75=> c0_n8_w75, 
            w76=> c0_n8_w76, 
            w77=> c0_n8_w77, 
            w78=> c0_n8_w78, 
            w79=> c0_n8_w79, 
            w80=> c0_n8_w80, 
            w81=> c0_n8_w81, 
            w82=> c0_n8_w82, 
            w83=> c0_n8_w83, 
            w84=> c0_n8_w84, 
            w85=> c0_n8_w85, 
            w86=> c0_n8_w86, 
            w87=> c0_n8_w87, 
            w88=> c0_n8_w88, 
            w89=> c0_n8_w89, 
            w90=> c0_n8_w90, 
            w91=> c0_n8_w91, 
            w92=> c0_n8_w92, 
            w93=> c0_n8_w93, 
            w94=> c0_n8_w94, 
            w95=> c0_n8_w95, 
            w96=> c0_n8_w96, 
            w97=> c0_n8_w97, 
            w98=> c0_n8_w98, 
            w99=> c0_n8_w99, 
            w100=> c0_n8_w100, 
            w101=> c0_n8_w101, 
            w102=> c0_n8_w102, 
            w103=> c0_n8_w103, 
            w104=> c0_n8_w104, 
            w105=> c0_n8_w105, 
            w106=> c0_n8_w106, 
            w107=> c0_n8_w107, 
            w108=> c0_n8_w108, 
            w109=> c0_n8_w109, 
            w110=> c0_n8_w110, 
            w111=> c0_n8_w111, 
            w112=> c0_n8_w112, 
            w113=> c0_n8_w113, 
            w114=> c0_n8_w114, 
            w115=> c0_n8_w115, 
            w116=> c0_n8_w116, 
            w117=> c0_n8_w117, 
            w118=> c0_n8_w118, 
            w119=> c0_n8_w119, 
            w120=> c0_n8_w120, 
            w121=> c0_n8_w121, 
            w122=> c0_n8_w122, 
            w123=> c0_n8_w123, 
            w124=> c0_n8_w124, 
            w125=> c0_n8_w125, 
            w126=> c0_n8_w126, 
            w127=> c0_n8_w127, 
            w128=> c0_n8_w128, 
            w129=> c0_n8_w129, 
            w130=> c0_n8_w130, 
            w131=> c0_n8_w131, 
            w132=> c0_n8_w132, 
            w133=> c0_n8_w133, 
            w134=> c0_n8_w134, 
            w135=> c0_n8_w135, 
            w136=> c0_n8_w136, 
            w137=> c0_n8_w137, 
            w138=> c0_n8_w138, 
            w139=> c0_n8_w139, 
            w140=> c0_n8_w140, 
            w141=> c0_n8_w141, 
            w142=> c0_n8_w142, 
            w143=> c0_n8_w143, 
            w144=> c0_n8_w144, 
            w145=> c0_n8_w145, 
            w146=> c0_n8_w146, 
            w147=> c0_n8_w147, 
            w148=> c0_n8_w148, 
            w149=> c0_n8_w149, 
            w150=> c0_n8_w150, 
            w151=> c0_n8_w151, 
            w152=> c0_n8_w152, 
            w153=> c0_n8_w153, 
            w154=> c0_n8_w154, 
            w155=> c0_n8_w155, 
            w156=> c0_n8_w156, 
            w157=> c0_n8_w157, 
            w158=> c0_n8_w158, 
            w159=> c0_n8_w159, 
            w160=> c0_n8_w160, 
            w161=> c0_n8_w161, 
            w162=> c0_n8_w162, 
            w163=> c0_n8_w163, 
            w164=> c0_n8_w164, 
            w165=> c0_n8_w165, 
            w166=> c0_n8_w166, 
            w167=> c0_n8_w167, 
            w168=> c0_n8_w168, 
            w169=> c0_n8_w169, 
            w170=> c0_n8_w170, 
            w171=> c0_n8_w171, 
            w172=> c0_n8_w172, 
            w173=> c0_n8_w173, 
            w174=> c0_n8_w174, 
            w175=> c0_n8_w175, 
            w176=> c0_n8_w176, 
            w177=> c0_n8_w177, 
            w178=> c0_n8_w178, 
            w179=> c0_n8_w179, 
            w180=> c0_n8_w180, 
            w181=> c0_n8_w181, 
            w182=> c0_n8_w182, 
            w183=> c0_n8_w183, 
            w184=> c0_n8_w184, 
            w185=> c0_n8_w185, 
            w186=> c0_n8_w186, 
            w187=> c0_n8_w187, 
            w188=> c0_n8_w188, 
            w189=> c0_n8_w189, 
            w190=> c0_n8_w190, 
            w191=> c0_n8_w191, 
            w192=> c0_n8_w192, 
            w193=> c0_n8_w193, 
            w194=> c0_n8_w194, 
            w195=> c0_n8_w195, 
            w196=> c0_n8_w196, 
            w197=> c0_n8_w197, 
            w198=> c0_n8_w198, 
            w199=> c0_n8_w199, 
            w200=> c0_n8_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n9_w1, 
            w2=> c0_n9_w2, 
            w3=> c0_n9_w3, 
            w4=> c0_n9_w4, 
            w5=> c0_n9_w5, 
            w6=> c0_n9_w6, 
            w7=> c0_n9_w7, 
            w8=> c0_n9_w8, 
            w9=> c0_n9_w9, 
            w10=> c0_n9_w10, 
            w11=> c0_n9_w11, 
            w12=> c0_n9_w12, 
            w13=> c0_n9_w13, 
            w14=> c0_n9_w14, 
            w15=> c0_n9_w15, 
            w16=> c0_n9_w16, 
            w17=> c0_n9_w17, 
            w18=> c0_n9_w18, 
            w19=> c0_n9_w19, 
            w20=> c0_n9_w20, 
            w21=> c0_n9_w21, 
            w22=> c0_n9_w22, 
            w23=> c0_n9_w23, 
            w24=> c0_n9_w24, 
            w25=> c0_n9_w25, 
            w26=> c0_n9_w26, 
            w27=> c0_n9_w27, 
            w28=> c0_n9_w28, 
            w29=> c0_n9_w29, 
            w30=> c0_n9_w30, 
            w31=> c0_n9_w31, 
            w32=> c0_n9_w32, 
            w33=> c0_n9_w33, 
            w34=> c0_n9_w34, 
            w35=> c0_n9_w35, 
            w36=> c0_n9_w36, 
            w37=> c0_n9_w37, 
            w38=> c0_n9_w38, 
            w39=> c0_n9_w39, 
            w40=> c0_n9_w40, 
            w41=> c0_n9_w41, 
            w42=> c0_n9_w42, 
            w43=> c0_n9_w43, 
            w44=> c0_n9_w44, 
            w45=> c0_n9_w45, 
            w46=> c0_n9_w46, 
            w47=> c0_n9_w47, 
            w48=> c0_n9_w48, 
            w49=> c0_n9_w49, 
            w50=> c0_n9_w50, 
            w51=> c0_n9_w51, 
            w52=> c0_n9_w52, 
            w53=> c0_n9_w53, 
            w54=> c0_n9_w54, 
            w55=> c0_n9_w55, 
            w56=> c0_n9_w56, 
            w57=> c0_n9_w57, 
            w58=> c0_n9_w58, 
            w59=> c0_n9_w59, 
            w60=> c0_n9_w60, 
            w61=> c0_n9_w61, 
            w62=> c0_n9_w62, 
            w63=> c0_n9_w63, 
            w64=> c0_n9_w64, 
            w65=> c0_n9_w65, 
            w66=> c0_n9_w66, 
            w67=> c0_n9_w67, 
            w68=> c0_n9_w68, 
            w69=> c0_n9_w69, 
            w70=> c0_n9_w70, 
            w71=> c0_n9_w71, 
            w72=> c0_n9_w72, 
            w73=> c0_n9_w73, 
            w74=> c0_n9_w74, 
            w75=> c0_n9_w75, 
            w76=> c0_n9_w76, 
            w77=> c0_n9_w77, 
            w78=> c0_n9_w78, 
            w79=> c0_n9_w79, 
            w80=> c0_n9_w80, 
            w81=> c0_n9_w81, 
            w82=> c0_n9_w82, 
            w83=> c0_n9_w83, 
            w84=> c0_n9_w84, 
            w85=> c0_n9_w85, 
            w86=> c0_n9_w86, 
            w87=> c0_n9_w87, 
            w88=> c0_n9_w88, 
            w89=> c0_n9_w89, 
            w90=> c0_n9_w90, 
            w91=> c0_n9_w91, 
            w92=> c0_n9_w92, 
            w93=> c0_n9_w93, 
            w94=> c0_n9_w94, 
            w95=> c0_n9_w95, 
            w96=> c0_n9_w96, 
            w97=> c0_n9_w97, 
            w98=> c0_n9_w98, 
            w99=> c0_n9_w99, 
            w100=> c0_n9_w100, 
            w101=> c0_n9_w101, 
            w102=> c0_n9_w102, 
            w103=> c0_n9_w103, 
            w104=> c0_n9_w104, 
            w105=> c0_n9_w105, 
            w106=> c0_n9_w106, 
            w107=> c0_n9_w107, 
            w108=> c0_n9_w108, 
            w109=> c0_n9_w109, 
            w110=> c0_n9_w110, 
            w111=> c0_n9_w111, 
            w112=> c0_n9_w112, 
            w113=> c0_n9_w113, 
            w114=> c0_n9_w114, 
            w115=> c0_n9_w115, 
            w116=> c0_n9_w116, 
            w117=> c0_n9_w117, 
            w118=> c0_n9_w118, 
            w119=> c0_n9_w119, 
            w120=> c0_n9_w120, 
            w121=> c0_n9_w121, 
            w122=> c0_n9_w122, 
            w123=> c0_n9_w123, 
            w124=> c0_n9_w124, 
            w125=> c0_n9_w125, 
            w126=> c0_n9_w126, 
            w127=> c0_n9_w127, 
            w128=> c0_n9_w128, 
            w129=> c0_n9_w129, 
            w130=> c0_n9_w130, 
            w131=> c0_n9_w131, 
            w132=> c0_n9_w132, 
            w133=> c0_n9_w133, 
            w134=> c0_n9_w134, 
            w135=> c0_n9_w135, 
            w136=> c0_n9_w136, 
            w137=> c0_n9_w137, 
            w138=> c0_n9_w138, 
            w139=> c0_n9_w139, 
            w140=> c0_n9_w140, 
            w141=> c0_n9_w141, 
            w142=> c0_n9_w142, 
            w143=> c0_n9_w143, 
            w144=> c0_n9_w144, 
            w145=> c0_n9_w145, 
            w146=> c0_n9_w146, 
            w147=> c0_n9_w147, 
            w148=> c0_n9_w148, 
            w149=> c0_n9_w149, 
            w150=> c0_n9_w150, 
            w151=> c0_n9_w151, 
            w152=> c0_n9_w152, 
            w153=> c0_n9_w153, 
            w154=> c0_n9_w154, 
            w155=> c0_n9_w155, 
            w156=> c0_n9_w156, 
            w157=> c0_n9_w157, 
            w158=> c0_n9_w158, 
            w159=> c0_n9_w159, 
            w160=> c0_n9_w160, 
            w161=> c0_n9_w161, 
            w162=> c0_n9_w162, 
            w163=> c0_n9_w163, 
            w164=> c0_n9_w164, 
            w165=> c0_n9_w165, 
            w166=> c0_n9_w166, 
            w167=> c0_n9_w167, 
            w168=> c0_n9_w168, 
            w169=> c0_n9_w169, 
            w170=> c0_n9_w170, 
            w171=> c0_n9_w171, 
            w172=> c0_n9_w172, 
            w173=> c0_n9_w173, 
            w174=> c0_n9_w174, 
            w175=> c0_n9_w175, 
            w176=> c0_n9_w176, 
            w177=> c0_n9_w177, 
            w178=> c0_n9_w178, 
            w179=> c0_n9_w179, 
            w180=> c0_n9_w180, 
            w181=> c0_n9_w181, 
            w182=> c0_n9_w182, 
            w183=> c0_n9_w183, 
            w184=> c0_n9_w184, 
            w185=> c0_n9_w185, 
            w186=> c0_n9_w186, 
            w187=> c0_n9_w187, 
            w188=> c0_n9_w188, 
            w189=> c0_n9_w189, 
            w190=> c0_n9_w190, 
            w191=> c0_n9_w191, 
            w192=> c0_n9_w192, 
            w193=> c0_n9_w193, 
            w194=> c0_n9_w194, 
            w195=> c0_n9_w195, 
            w196=> c0_n9_w196, 
            w197=> c0_n9_w197, 
            w198=> c0_n9_w198, 
            w199=> c0_n9_w199, 
            w200=> c0_n9_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n9_y
   );           
            
neuron_inst_10: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n10_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n10_w1, 
            w2=> c0_n10_w2, 
            w3=> c0_n10_w3, 
            w4=> c0_n10_w4, 
            w5=> c0_n10_w5, 
            w6=> c0_n10_w6, 
            w7=> c0_n10_w7, 
            w8=> c0_n10_w8, 
            w9=> c0_n10_w9, 
            w10=> c0_n10_w10, 
            w11=> c0_n10_w11, 
            w12=> c0_n10_w12, 
            w13=> c0_n10_w13, 
            w14=> c0_n10_w14, 
            w15=> c0_n10_w15, 
            w16=> c0_n10_w16, 
            w17=> c0_n10_w17, 
            w18=> c0_n10_w18, 
            w19=> c0_n10_w19, 
            w20=> c0_n10_w20, 
            w21=> c0_n10_w21, 
            w22=> c0_n10_w22, 
            w23=> c0_n10_w23, 
            w24=> c0_n10_w24, 
            w25=> c0_n10_w25, 
            w26=> c0_n10_w26, 
            w27=> c0_n10_w27, 
            w28=> c0_n10_w28, 
            w29=> c0_n10_w29, 
            w30=> c0_n10_w30, 
            w31=> c0_n10_w31, 
            w32=> c0_n10_w32, 
            w33=> c0_n10_w33, 
            w34=> c0_n10_w34, 
            w35=> c0_n10_w35, 
            w36=> c0_n10_w36, 
            w37=> c0_n10_w37, 
            w38=> c0_n10_w38, 
            w39=> c0_n10_w39, 
            w40=> c0_n10_w40, 
            w41=> c0_n10_w41, 
            w42=> c0_n10_w42, 
            w43=> c0_n10_w43, 
            w44=> c0_n10_w44, 
            w45=> c0_n10_w45, 
            w46=> c0_n10_w46, 
            w47=> c0_n10_w47, 
            w48=> c0_n10_w48, 
            w49=> c0_n10_w49, 
            w50=> c0_n10_w50, 
            w51=> c0_n10_w51, 
            w52=> c0_n10_w52, 
            w53=> c0_n10_w53, 
            w54=> c0_n10_w54, 
            w55=> c0_n10_w55, 
            w56=> c0_n10_w56, 
            w57=> c0_n10_w57, 
            w58=> c0_n10_w58, 
            w59=> c0_n10_w59, 
            w60=> c0_n10_w60, 
            w61=> c0_n10_w61, 
            w62=> c0_n10_w62, 
            w63=> c0_n10_w63, 
            w64=> c0_n10_w64, 
            w65=> c0_n10_w65, 
            w66=> c0_n10_w66, 
            w67=> c0_n10_w67, 
            w68=> c0_n10_w68, 
            w69=> c0_n10_w69, 
            w70=> c0_n10_w70, 
            w71=> c0_n10_w71, 
            w72=> c0_n10_w72, 
            w73=> c0_n10_w73, 
            w74=> c0_n10_w74, 
            w75=> c0_n10_w75, 
            w76=> c0_n10_w76, 
            w77=> c0_n10_w77, 
            w78=> c0_n10_w78, 
            w79=> c0_n10_w79, 
            w80=> c0_n10_w80, 
            w81=> c0_n10_w81, 
            w82=> c0_n10_w82, 
            w83=> c0_n10_w83, 
            w84=> c0_n10_w84, 
            w85=> c0_n10_w85, 
            w86=> c0_n10_w86, 
            w87=> c0_n10_w87, 
            w88=> c0_n10_w88, 
            w89=> c0_n10_w89, 
            w90=> c0_n10_w90, 
            w91=> c0_n10_w91, 
            w92=> c0_n10_w92, 
            w93=> c0_n10_w93, 
            w94=> c0_n10_w94, 
            w95=> c0_n10_w95, 
            w96=> c0_n10_w96, 
            w97=> c0_n10_w97, 
            w98=> c0_n10_w98, 
            w99=> c0_n10_w99, 
            w100=> c0_n10_w100, 
            w101=> c0_n10_w101, 
            w102=> c0_n10_w102, 
            w103=> c0_n10_w103, 
            w104=> c0_n10_w104, 
            w105=> c0_n10_w105, 
            w106=> c0_n10_w106, 
            w107=> c0_n10_w107, 
            w108=> c0_n10_w108, 
            w109=> c0_n10_w109, 
            w110=> c0_n10_w110, 
            w111=> c0_n10_w111, 
            w112=> c0_n10_w112, 
            w113=> c0_n10_w113, 
            w114=> c0_n10_w114, 
            w115=> c0_n10_w115, 
            w116=> c0_n10_w116, 
            w117=> c0_n10_w117, 
            w118=> c0_n10_w118, 
            w119=> c0_n10_w119, 
            w120=> c0_n10_w120, 
            w121=> c0_n10_w121, 
            w122=> c0_n10_w122, 
            w123=> c0_n10_w123, 
            w124=> c0_n10_w124, 
            w125=> c0_n10_w125, 
            w126=> c0_n10_w126, 
            w127=> c0_n10_w127, 
            w128=> c0_n10_w128, 
            w129=> c0_n10_w129, 
            w130=> c0_n10_w130, 
            w131=> c0_n10_w131, 
            w132=> c0_n10_w132, 
            w133=> c0_n10_w133, 
            w134=> c0_n10_w134, 
            w135=> c0_n10_w135, 
            w136=> c0_n10_w136, 
            w137=> c0_n10_w137, 
            w138=> c0_n10_w138, 
            w139=> c0_n10_w139, 
            w140=> c0_n10_w140, 
            w141=> c0_n10_w141, 
            w142=> c0_n10_w142, 
            w143=> c0_n10_w143, 
            w144=> c0_n10_w144, 
            w145=> c0_n10_w145, 
            w146=> c0_n10_w146, 
            w147=> c0_n10_w147, 
            w148=> c0_n10_w148, 
            w149=> c0_n10_w149, 
            w150=> c0_n10_w150, 
            w151=> c0_n10_w151, 
            w152=> c0_n10_w152, 
            w153=> c0_n10_w153, 
            w154=> c0_n10_w154, 
            w155=> c0_n10_w155, 
            w156=> c0_n10_w156, 
            w157=> c0_n10_w157, 
            w158=> c0_n10_w158, 
            w159=> c0_n10_w159, 
            w160=> c0_n10_w160, 
            w161=> c0_n10_w161, 
            w162=> c0_n10_w162, 
            w163=> c0_n10_w163, 
            w164=> c0_n10_w164, 
            w165=> c0_n10_w165, 
            w166=> c0_n10_w166, 
            w167=> c0_n10_w167, 
            w168=> c0_n10_w168, 
            w169=> c0_n10_w169, 
            w170=> c0_n10_w170, 
            w171=> c0_n10_w171, 
            w172=> c0_n10_w172, 
            w173=> c0_n10_w173, 
            w174=> c0_n10_w174, 
            w175=> c0_n10_w175, 
            w176=> c0_n10_w176, 
            w177=> c0_n10_w177, 
            w178=> c0_n10_w178, 
            w179=> c0_n10_w179, 
            w180=> c0_n10_w180, 
            w181=> c0_n10_w181, 
            w182=> c0_n10_w182, 
            w183=> c0_n10_w183, 
            w184=> c0_n10_w184, 
            w185=> c0_n10_w185, 
            w186=> c0_n10_w186, 
            w187=> c0_n10_w187, 
            w188=> c0_n10_w188, 
            w189=> c0_n10_w189, 
            w190=> c0_n10_w190, 
            w191=> c0_n10_w191, 
            w192=> c0_n10_w192, 
            w193=> c0_n10_w193, 
            w194=> c0_n10_w194, 
            w195=> c0_n10_w195, 
            w196=> c0_n10_w196, 
            w197=> c0_n10_w197, 
            w198=> c0_n10_w198, 
            w199=> c0_n10_w199, 
            w200=> c0_n10_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n10_y
   );           
            
neuron_inst_11: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n11_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n11_w1, 
            w2=> c0_n11_w2, 
            w3=> c0_n11_w3, 
            w4=> c0_n11_w4, 
            w5=> c0_n11_w5, 
            w6=> c0_n11_w6, 
            w7=> c0_n11_w7, 
            w8=> c0_n11_w8, 
            w9=> c0_n11_w9, 
            w10=> c0_n11_w10, 
            w11=> c0_n11_w11, 
            w12=> c0_n11_w12, 
            w13=> c0_n11_w13, 
            w14=> c0_n11_w14, 
            w15=> c0_n11_w15, 
            w16=> c0_n11_w16, 
            w17=> c0_n11_w17, 
            w18=> c0_n11_w18, 
            w19=> c0_n11_w19, 
            w20=> c0_n11_w20, 
            w21=> c0_n11_w21, 
            w22=> c0_n11_w22, 
            w23=> c0_n11_w23, 
            w24=> c0_n11_w24, 
            w25=> c0_n11_w25, 
            w26=> c0_n11_w26, 
            w27=> c0_n11_w27, 
            w28=> c0_n11_w28, 
            w29=> c0_n11_w29, 
            w30=> c0_n11_w30, 
            w31=> c0_n11_w31, 
            w32=> c0_n11_w32, 
            w33=> c0_n11_w33, 
            w34=> c0_n11_w34, 
            w35=> c0_n11_w35, 
            w36=> c0_n11_w36, 
            w37=> c0_n11_w37, 
            w38=> c0_n11_w38, 
            w39=> c0_n11_w39, 
            w40=> c0_n11_w40, 
            w41=> c0_n11_w41, 
            w42=> c0_n11_w42, 
            w43=> c0_n11_w43, 
            w44=> c0_n11_w44, 
            w45=> c0_n11_w45, 
            w46=> c0_n11_w46, 
            w47=> c0_n11_w47, 
            w48=> c0_n11_w48, 
            w49=> c0_n11_w49, 
            w50=> c0_n11_w50, 
            w51=> c0_n11_w51, 
            w52=> c0_n11_w52, 
            w53=> c0_n11_w53, 
            w54=> c0_n11_w54, 
            w55=> c0_n11_w55, 
            w56=> c0_n11_w56, 
            w57=> c0_n11_w57, 
            w58=> c0_n11_w58, 
            w59=> c0_n11_w59, 
            w60=> c0_n11_w60, 
            w61=> c0_n11_w61, 
            w62=> c0_n11_w62, 
            w63=> c0_n11_w63, 
            w64=> c0_n11_w64, 
            w65=> c0_n11_w65, 
            w66=> c0_n11_w66, 
            w67=> c0_n11_w67, 
            w68=> c0_n11_w68, 
            w69=> c0_n11_w69, 
            w70=> c0_n11_w70, 
            w71=> c0_n11_w71, 
            w72=> c0_n11_w72, 
            w73=> c0_n11_w73, 
            w74=> c0_n11_w74, 
            w75=> c0_n11_w75, 
            w76=> c0_n11_w76, 
            w77=> c0_n11_w77, 
            w78=> c0_n11_w78, 
            w79=> c0_n11_w79, 
            w80=> c0_n11_w80, 
            w81=> c0_n11_w81, 
            w82=> c0_n11_w82, 
            w83=> c0_n11_w83, 
            w84=> c0_n11_w84, 
            w85=> c0_n11_w85, 
            w86=> c0_n11_w86, 
            w87=> c0_n11_w87, 
            w88=> c0_n11_w88, 
            w89=> c0_n11_w89, 
            w90=> c0_n11_w90, 
            w91=> c0_n11_w91, 
            w92=> c0_n11_w92, 
            w93=> c0_n11_w93, 
            w94=> c0_n11_w94, 
            w95=> c0_n11_w95, 
            w96=> c0_n11_w96, 
            w97=> c0_n11_w97, 
            w98=> c0_n11_w98, 
            w99=> c0_n11_w99, 
            w100=> c0_n11_w100, 
            w101=> c0_n11_w101, 
            w102=> c0_n11_w102, 
            w103=> c0_n11_w103, 
            w104=> c0_n11_w104, 
            w105=> c0_n11_w105, 
            w106=> c0_n11_w106, 
            w107=> c0_n11_w107, 
            w108=> c0_n11_w108, 
            w109=> c0_n11_w109, 
            w110=> c0_n11_w110, 
            w111=> c0_n11_w111, 
            w112=> c0_n11_w112, 
            w113=> c0_n11_w113, 
            w114=> c0_n11_w114, 
            w115=> c0_n11_w115, 
            w116=> c0_n11_w116, 
            w117=> c0_n11_w117, 
            w118=> c0_n11_w118, 
            w119=> c0_n11_w119, 
            w120=> c0_n11_w120, 
            w121=> c0_n11_w121, 
            w122=> c0_n11_w122, 
            w123=> c0_n11_w123, 
            w124=> c0_n11_w124, 
            w125=> c0_n11_w125, 
            w126=> c0_n11_w126, 
            w127=> c0_n11_w127, 
            w128=> c0_n11_w128, 
            w129=> c0_n11_w129, 
            w130=> c0_n11_w130, 
            w131=> c0_n11_w131, 
            w132=> c0_n11_w132, 
            w133=> c0_n11_w133, 
            w134=> c0_n11_w134, 
            w135=> c0_n11_w135, 
            w136=> c0_n11_w136, 
            w137=> c0_n11_w137, 
            w138=> c0_n11_w138, 
            w139=> c0_n11_w139, 
            w140=> c0_n11_w140, 
            w141=> c0_n11_w141, 
            w142=> c0_n11_w142, 
            w143=> c0_n11_w143, 
            w144=> c0_n11_w144, 
            w145=> c0_n11_w145, 
            w146=> c0_n11_w146, 
            w147=> c0_n11_w147, 
            w148=> c0_n11_w148, 
            w149=> c0_n11_w149, 
            w150=> c0_n11_w150, 
            w151=> c0_n11_w151, 
            w152=> c0_n11_w152, 
            w153=> c0_n11_w153, 
            w154=> c0_n11_w154, 
            w155=> c0_n11_w155, 
            w156=> c0_n11_w156, 
            w157=> c0_n11_w157, 
            w158=> c0_n11_w158, 
            w159=> c0_n11_w159, 
            w160=> c0_n11_w160, 
            w161=> c0_n11_w161, 
            w162=> c0_n11_w162, 
            w163=> c0_n11_w163, 
            w164=> c0_n11_w164, 
            w165=> c0_n11_w165, 
            w166=> c0_n11_w166, 
            w167=> c0_n11_w167, 
            w168=> c0_n11_w168, 
            w169=> c0_n11_w169, 
            w170=> c0_n11_w170, 
            w171=> c0_n11_w171, 
            w172=> c0_n11_w172, 
            w173=> c0_n11_w173, 
            w174=> c0_n11_w174, 
            w175=> c0_n11_w175, 
            w176=> c0_n11_w176, 
            w177=> c0_n11_w177, 
            w178=> c0_n11_w178, 
            w179=> c0_n11_w179, 
            w180=> c0_n11_w180, 
            w181=> c0_n11_w181, 
            w182=> c0_n11_w182, 
            w183=> c0_n11_w183, 
            w184=> c0_n11_w184, 
            w185=> c0_n11_w185, 
            w186=> c0_n11_w186, 
            w187=> c0_n11_w187, 
            w188=> c0_n11_w188, 
            w189=> c0_n11_w189, 
            w190=> c0_n11_w190, 
            w191=> c0_n11_w191, 
            w192=> c0_n11_w192, 
            w193=> c0_n11_w193, 
            w194=> c0_n11_w194, 
            w195=> c0_n11_w195, 
            w196=> c0_n11_w196, 
            w197=> c0_n11_w197, 
            w198=> c0_n11_w198, 
            w199=> c0_n11_w199, 
            w200=> c0_n11_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n11_y
   );           
            
neuron_inst_12: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n12_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n12_w1, 
            w2=> c0_n12_w2, 
            w3=> c0_n12_w3, 
            w4=> c0_n12_w4, 
            w5=> c0_n12_w5, 
            w6=> c0_n12_w6, 
            w7=> c0_n12_w7, 
            w8=> c0_n12_w8, 
            w9=> c0_n12_w9, 
            w10=> c0_n12_w10, 
            w11=> c0_n12_w11, 
            w12=> c0_n12_w12, 
            w13=> c0_n12_w13, 
            w14=> c0_n12_w14, 
            w15=> c0_n12_w15, 
            w16=> c0_n12_w16, 
            w17=> c0_n12_w17, 
            w18=> c0_n12_w18, 
            w19=> c0_n12_w19, 
            w20=> c0_n12_w20, 
            w21=> c0_n12_w21, 
            w22=> c0_n12_w22, 
            w23=> c0_n12_w23, 
            w24=> c0_n12_w24, 
            w25=> c0_n12_w25, 
            w26=> c0_n12_w26, 
            w27=> c0_n12_w27, 
            w28=> c0_n12_w28, 
            w29=> c0_n12_w29, 
            w30=> c0_n12_w30, 
            w31=> c0_n12_w31, 
            w32=> c0_n12_w32, 
            w33=> c0_n12_w33, 
            w34=> c0_n12_w34, 
            w35=> c0_n12_w35, 
            w36=> c0_n12_w36, 
            w37=> c0_n12_w37, 
            w38=> c0_n12_w38, 
            w39=> c0_n12_w39, 
            w40=> c0_n12_w40, 
            w41=> c0_n12_w41, 
            w42=> c0_n12_w42, 
            w43=> c0_n12_w43, 
            w44=> c0_n12_w44, 
            w45=> c0_n12_w45, 
            w46=> c0_n12_w46, 
            w47=> c0_n12_w47, 
            w48=> c0_n12_w48, 
            w49=> c0_n12_w49, 
            w50=> c0_n12_w50, 
            w51=> c0_n12_w51, 
            w52=> c0_n12_w52, 
            w53=> c0_n12_w53, 
            w54=> c0_n12_w54, 
            w55=> c0_n12_w55, 
            w56=> c0_n12_w56, 
            w57=> c0_n12_w57, 
            w58=> c0_n12_w58, 
            w59=> c0_n12_w59, 
            w60=> c0_n12_w60, 
            w61=> c0_n12_w61, 
            w62=> c0_n12_w62, 
            w63=> c0_n12_w63, 
            w64=> c0_n12_w64, 
            w65=> c0_n12_w65, 
            w66=> c0_n12_w66, 
            w67=> c0_n12_w67, 
            w68=> c0_n12_w68, 
            w69=> c0_n12_w69, 
            w70=> c0_n12_w70, 
            w71=> c0_n12_w71, 
            w72=> c0_n12_w72, 
            w73=> c0_n12_w73, 
            w74=> c0_n12_w74, 
            w75=> c0_n12_w75, 
            w76=> c0_n12_w76, 
            w77=> c0_n12_w77, 
            w78=> c0_n12_w78, 
            w79=> c0_n12_w79, 
            w80=> c0_n12_w80, 
            w81=> c0_n12_w81, 
            w82=> c0_n12_w82, 
            w83=> c0_n12_w83, 
            w84=> c0_n12_w84, 
            w85=> c0_n12_w85, 
            w86=> c0_n12_w86, 
            w87=> c0_n12_w87, 
            w88=> c0_n12_w88, 
            w89=> c0_n12_w89, 
            w90=> c0_n12_w90, 
            w91=> c0_n12_w91, 
            w92=> c0_n12_w92, 
            w93=> c0_n12_w93, 
            w94=> c0_n12_w94, 
            w95=> c0_n12_w95, 
            w96=> c0_n12_w96, 
            w97=> c0_n12_w97, 
            w98=> c0_n12_w98, 
            w99=> c0_n12_w99, 
            w100=> c0_n12_w100, 
            w101=> c0_n12_w101, 
            w102=> c0_n12_w102, 
            w103=> c0_n12_w103, 
            w104=> c0_n12_w104, 
            w105=> c0_n12_w105, 
            w106=> c0_n12_w106, 
            w107=> c0_n12_w107, 
            w108=> c0_n12_w108, 
            w109=> c0_n12_w109, 
            w110=> c0_n12_w110, 
            w111=> c0_n12_w111, 
            w112=> c0_n12_w112, 
            w113=> c0_n12_w113, 
            w114=> c0_n12_w114, 
            w115=> c0_n12_w115, 
            w116=> c0_n12_w116, 
            w117=> c0_n12_w117, 
            w118=> c0_n12_w118, 
            w119=> c0_n12_w119, 
            w120=> c0_n12_w120, 
            w121=> c0_n12_w121, 
            w122=> c0_n12_w122, 
            w123=> c0_n12_w123, 
            w124=> c0_n12_w124, 
            w125=> c0_n12_w125, 
            w126=> c0_n12_w126, 
            w127=> c0_n12_w127, 
            w128=> c0_n12_w128, 
            w129=> c0_n12_w129, 
            w130=> c0_n12_w130, 
            w131=> c0_n12_w131, 
            w132=> c0_n12_w132, 
            w133=> c0_n12_w133, 
            w134=> c0_n12_w134, 
            w135=> c0_n12_w135, 
            w136=> c0_n12_w136, 
            w137=> c0_n12_w137, 
            w138=> c0_n12_w138, 
            w139=> c0_n12_w139, 
            w140=> c0_n12_w140, 
            w141=> c0_n12_w141, 
            w142=> c0_n12_w142, 
            w143=> c0_n12_w143, 
            w144=> c0_n12_w144, 
            w145=> c0_n12_w145, 
            w146=> c0_n12_w146, 
            w147=> c0_n12_w147, 
            w148=> c0_n12_w148, 
            w149=> c0_n12_w149, 
            w150=> c0_n12_w150, 
            w151=> c0_n12_w151, 
            w152=> c0_n12_w152, 
            w153=> c0_n12_w153, 
            w154=> c0_n12_w154, 
            w155=> c0_n12_w155, 
            w156=> c0_n12_w156, 
            w157=> c0_n12_w157, 
            w158=> c0_n12_w158, 
            w159=> c0_n12_w159, 
            w160=> c0_n12_w160, 
            w161=> c0_n12_w161, 
            w162=> c0_n12_w162, 
            w163=> c0_n12_w163, 
            w164=> c0_n12_w164, 
            w165=> c0_n12_w165, 
            w166=> c0_n12_w166, 
            w167=> c0_n12_w167, 
            w168=> c0_n12_w168, 
            w169=> c0_n12_w169, 
            w170=> c0_n12_w170, 
            w171=> c0_n12_w171, 
            w172=> c0_n12_w172, 
            w173=> c0_n12_w173, 
            w174=> c0_n12_w174, 
            w175=> c0_n12_w175, 
            w176=> c0_n12_w176, 
            w177=> c0_n12_w177, 
            w178=> c0_n12_w178, 
            w179=> c0_n12_w179, 
            w180=> c0_n12_w180, 
            w181=> c0_n12_w181, 
            w182=> c0_n12_w182, 
            w183=> c0_n12_w183, 
            w184=> c0_n12_w184, 
            w185=> c0_n12_w185, 
            w186=> c0_n12_w186, 
            w187=> c0_n12_w187, 
            w188=> c0_n12_w188, 
            w189=> c0_n12_w189, 
            w190=> c0_n12_w190, 
            w191=> c0_n12_w191, 
            w192=> c0_n12_w192, 
            w193=> c0_n12_w193, 
            w194=> c0_n12_w194, 
            w195=> c0_n12_w195, 
            w196=> c0_n12_w196, 
            w197=> c0_n12_w197, 
            w198=> c0_n12_w198, 
            w199=> c0_n12_w199, 
            w200=> c0_n12_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n12_y
   );           
            
neuron_inst_13: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n13_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n13_w1, 
            w2=> c0_n13_w2, 
            w3=> c0_n13_w3, 
            w4=> c0_n13_w4, 
            w5=> c0_n13_w5, 
            w6=> c0_n13_w6, 
            w7=> c0_n13_w7, 
            w8=> c0_n13_w8, 
            w9=> c0_n13_w9, 
            w10=> c0_n13_w10, 
            w11=> c0_n13_w11, 
            w12=> c0_n13_w12, 
            w13=> c0_n13_w13, 
            w14=> c0_n13_w14, 
            w15=> c0_n13_w15, 
            w16=> c0_n13_w16, 
            w17=> c0_n13_w17, 
            w18=> c0_n13_w18, 
            w19=> c0_n13_w19, 
            w20=> c0_n13_w20, 
            w21=> c0_n13_w21, 
            w22=> c0_n13_w22, 
            w23=> c0_n13_w23, 
            w24=> c0_n13_w24, 
            w25=> c0_n13_w25, 
            w26=> c0_n13_w26, 
            w27=> c0_n13_w27, 
            w28=> c0_n13_w28, 
            w29=> c0_n13_w29, 
            w30=> c0_n13_w30, 
            w31=> c0_n13_w31, 
            w32=> c0_n13_w32, 
            w33=> c0_n13_w33, 
            w34=> c0_n13_w34, 
            w35=> c0_n13_w35, 
            w36=> c0_n13_w36, 
            w37=> c0_n13_w37, 
            w38=> c0_n13_w38, 
            w39=> c0_n13_w39, 
            w40=> c0_n13_w40, 
            w41=> c0_n13_w41, 
            w42=> c0_n13_w42, 
            w43=> c0_n13_w43, 
            w44=> c0_n13_w44, 
            w45=> c0_n13_w45, 
            w46=> c0_n13_w46, 
            w47=> c0_n13_w47, 
            w48=> c0_n13_w48, 
            w49=> c0_n13_w49, 
            w50=> c0_n13_w50, 
            w51=> c0_n13_w51, 
            w52=> c0_n13_w52, 
            w53=> c0_n13_w53, 
            w54=> c0_n13_w54, 
            w55=> c0_n13_w55, 
            w56=> c0_n13_w56, 
            w57=> c0_n13_w57, 
            w58=> c0_n13_w58, 
            w59=> c0_n13_w59, 
            w60=> c0_n13_w60, 
            w61=> c0_n13_w61, 
            w62=> c0_n13_w62, 
            w63=> c0_n13_w63, 
            w64=> c0_n13_w64, 
            w65=> c0_n13_w65, 
            w66=> c0_n13_w66, 
            w67=> c0_n13_w67, 
            w68=> c0_n13_w68, 
            w69=> c0_n13_w69, 
            w70=> c0_n13_w70, 
            w71=> c0_n13_w71, 
            w72=> c0_n13_w72, 
            w73=> c0_n13_w73, 
            w74=> c0_n13_w74, 
            w75=> c0_n13_w75, 
            w76=> c0_n13_w76, 
            w77=> c0_n13_w77, 
            w78=> c0_n13_w78, 
            w79=> c0_n13_w79, 
            w80=> c0_n13_w80, 
            w81=> c0_n13_w81, 
            w82=> c0_n13_w82, 
            w83=> c0_n13_w83, 
            w84=> c0_n13_w84, 
            w85=> c0_n13_w85, 
            w86=> c0_n13_w86, 
            w87=> c0_n13_w87, 
            w88=> c0_n13_w88, 
            w89=> c0_n13_w89, 
            w90=> c0_n13_w90, 
            w91=> c0_n13_w91, 
            w92=> c0_n13_w92, 
            w93=> c0_n13_w93, 
            w94=> c0_n13_w94, 
            w95=> c0_n13_w95, 
            w96=> c0_n13_w96, 
            w97=> c0_n13_w97, 
            w98=> c0_n13_w98, 
            w99=> c0_n13_w99, 
            w100=> c0_n13_w100, 
            w101=> c0_n13_w101, 
            w102=> c0_n13_w102, 
            w103=> c0_n13_w103, 
            w104=> c0_n13_w104, 
            w105=> c0_n13_w105, 
            w106=> c0_n13_w106, 
            w107=> c0_n13_w107, 
            w108=> c0_n13_w108, 
            w109=> c0_n13_w109, 
            w110=> c0_n13_w110, 
            w111=> c0_n13_w111, 
            w112=> c0_n13_w112, 
            w113=> c0_n13_w113, 
            w114=> c0_n13_w114, 
            w115=> c0_n13_w115, 
            w116=> c0_n13_w116, 
            w117=> c0_n13_w117, 
            w118=> c0_n13_w118, 
            w119=> c0_n13_w119, 
            w120=> c0_n13_w120, 
            w121=> c0_n13_w121, 
            w122=> c0_n13_w122, 
            w123=> c0_n13_w123, 
            w124=> c0_n13_w124, 
            w125=> c0_n13_w125, 
            w126=> c0_n13_w126, 
            w127=> c0_n13_w127, 
            w128=> c0_n13_w128, 
            w129=> c0_n13_w129, 
            w130=> c0_n13_w130, 
            w131=> c0_n13_w131, 
            w132=> c0_n13_w132, 
            w133=> c0_n13_w133, 
            w134=> c0_n13_w134, 
            w135=> c0_n13_w135, 
            w136=> c0_n13_w136, 
            w137=> c0_n13_w137, 
            w138=> c0_n13_w138, 
            w139=> c0_n13_w139, 
            w140=> c0_n13_w140, 
            w141=> c0_n13_w141, 
            w142=> c0_n13_w142, 
            w143=> c0_n13_w143, 
            w144=> c0_n13_w144, 
            w145=> c0_n13_w145, 
            w146=> c0_n13_w146, 
            w147=> c0_n13_w147, 
            w148=> c0_n13_w148, 
            w149=> c0_n13_w149, 
            w150=> c0_n13_w150, 
            w151=> c0_n13_w151, 
            w152=> c0_n13_w152, 
            w153=> c0_n13_w153, 
            w154=> c0_n13_w154, 
            w155=> c0_n13_w155, 
            w156=> c0_n13_w156, 
            w157=> c0_n13_w157, 
            w158=> c0_n13_w158, 
            w159=> c0_n13_w159, 
            w160=> c0_n13_w160, 
            w161=> c0_n13_w161, 
            w162=> c0_n13_w162, 
            w163=> c0_n13_w163, 
            w164=> c0_n13_w164, 
            w165=> c0_n13_w165, 
            w166=> c0_n13_w166, 
            w167=> c0_n13_w167, 
            w168=> c0_n13_w168, 
            w169=> c0_n13_w169, 
            w170=> c0_n13_w170, 
            w171=> c0_n13_w171, 
            w172=> c0_n13_w172, 
            w173=> c0_n13_w173, 
            w174=> c0_n13_w174, 
            w175=> c0_n13_w175, 
            w176=> c0_n13_w176, 
            w177=> c0_n13_w177, 
            w178=> c0_n13_w178, 
            w179=> c0_n13_w179, 
            w180=> c0_n13_w180, 
            w181=> c0_n13_w181, 
            w182=> c0_n13_w182, 
            w183=> c0_n13_w183, 
            w184=> c0_n13_w184, 
            w185=> c0_n13_w185, 
            w186=> c0_n13_w186, 
            w187=> c0_n13_w187, 
            w188=> c0_n13_w188, 
            w189=> c0_n13_w189, 
            w190=> c0_n13_w190, 
            w191=> c0_n13_w191, 
            w192=> c0_n13_w192, 
            w193=> c0_n13_w193, 
            w194=> c0_n13_w194, 
            w195=> c0_n13_w195, 
            w196=> c0_n13_w196, 
            w197=> c0_n13_w197, 
            w198=> c0_n13_w198, 
            w199=> c0_n13_w199, 
            w200=> c0_n13_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n13_y
   );           
            
neuron_inst_14: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n14_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n14_w1, 
            w2=> c0_n14_w2, 
            w3=> c0_n14_w3, 
            w4=> c0_n14_w4, 
            w5=> c0_n14_w5, 
            w6=> c0_n14_w6, 
            w7=> c0_n14_w7, 
            w8=> c0_n14_w8, 
            w9=> c0_n14_w9, 
            w10=> c0_n14_w10, 
            w11=> c0_n14_w11, 
            w12=> c0_n14_w12, 
            w13=> c0_n14_w13, 
            w14=> c0_n14_w14, 
            w15=> c0_n14_w15, 
            w16=> c0_n14_w16, 
            w17=> c0_n14_w17, 
            w18=> c0_n14_w18, 
            w19=> c0_n14_w19, 
            w20=> c0_n14_w20, 
            w21=> c0_n14_w21, 
            w22=> c0_n14_w22, 
            w23=> c0_n14_w23, 
            w24=> c0_n14_w24, 
            w25=> c0_n14_w25, 
            w26=> c0_n14_w26, 
            w27=> c0_n14_w27, 
            w28=> c0_n14_w28, 
            w29=> c0_n14_w29, 
            w30=> c0_n14_w30, 
            w31=> c0_n14_w31, 
            w32=> c0_n14_w32, 
            w33=> c0_n14_w33, 
            w34=> c0_n14_w34, 
            w35=> c0_n14_w35, 
            w36=> c0_n14_w36, 
            w37=> c0_n14_w37, 
            w38=> c0_n14_w38, 
            w39=> c0_n14_w39, 
            w40=> c0_n14_w40, 
            w41=> c0_n14_w41, 
            w42=> c0_n14_w42, 
            w43=> c0_n14_w43, 
            w44=> c0_n14_w44, 
            w45=> c0_n14_w45, 
            w46=> c0_n14_w46, 
            w47=> c0_n14_w47, 
            w48=> c0_n14_w48, 
            w49=> c0_n14_w49, 
            w50=> c0_n14_w50, 
            w51=> c0_n14_w51, 
            w52=> c0_n14_w52, 
            w53=> c0_n14_w53, 
            w54=> c0_n14_w54, 
            w55=> c0_n14_w55, 
            w56=> c0_n14_w56, 
            w57=> c0_n14_w57, 
            w58=> c0_n14_w58, 
            w59=> c0_n14_w59, 
            w60=> c0_n14_w60, 
            w61=> c0_n14_w61, 
            w62=> c0_n14_w62, 
            w63=> c0_n14_w63, 
            w64=> c0_n14_w64, 
            w65=> c0_n14_w65, 
            w66=> c0_n14_w66, 
            w67=> c0_n14_w67, 
            w68=> c0_n14_w68, 
            w69=> c0_n14_w69, 
            w70=> c0_n14_w70, 
            w71=> c0_n14_w71, 
            w72=> c0_n14_w72, 
            w73=> c0_n14_w73, 
            w74=> c0_n14_w74, 
            w75=> c0_n14_w75, 
            w76=> c0_n14_w76, 
            w77=> c0_n14_w77, 
            w78=> c0_n14_w78, 
            w79=> c0_n14_w79, 
            w80=> c0_n14_w80, 
            w81=> c0_n14_w81, 
            w82=> c0_n14_w82, 
            w83=> c0_n14_w83, 
            w84=> c0_n14_w84, 
            w85=> c0_n14_w85, 
            w86=> c0_n14_w86, 
            w87=> c0_n14_w87, 
            w88=> c0_n14_w88, 
            w89=> c0_n14_w89, 
            w90=> c0_n14_w90, 
            w91=> c0_n14_w91, 
            w92=> c0_n14_w92, 
            w93=> c0_n14_w93, 
            w94=> c0_n14_w94, 
            w95=> c0_n14_w95, 
            w96=> c0_n14_w96, 
            w97=> c0_n14_w97, 
            w98=> c0_n14_w98, 
            w99=> c0_n14_w99, 
            w100=> c0_n14_w100, 
            w101=> c0_n14_w101, 
            w102=> c0_n14_w102, 
            w103=> c0_n14_w103, 
            w104=> c0_n14_w104, 
            w105=> c0_n14_w105, 
            w106=> c0_n14_w106, 
            w107=> c0_n14_w107, 
            w108=> c0_n14_w108, 
            w109=> c0_n14_w109, 
            w110=> c0_n14_w110, 
            w111=> c0_n14_w111, 
            w112=> c0_n14_w112, 
            w113=> c0_n14_w113, 
            w114=> c0_n14_w114, 
            w115=> c0_n14_w115, 
            w116=> c0_n14_w116, 
            w117=> c0_n14_w117, 
            w118=> c0_n14_w118, 
            w119=> c0_n14_w119, 
            w120=> c0_n14_w120, 
            w121=> c0_n14_w121, 
            w122=> c0_n14_w122, 
            w123=> c0_n14_w123, 
            w124=> c0_n14_w124, 
            w125=> c0_n14_w125, 
            w126=> c0_n14_w126, 
            w127=> c0_n14_w127, 
            w128=> c0_n14_w128, 
            w129=> c0_n14_w129, 
            w130=> c0_n14_w130, 
            w131=> c0_n14_w131, 
            w132=> c0_n14_w132, 
            w133=> c0_n14_w133, 
            w134=> c0_n14_w134, 
            w135=> c0_n14_w135, 
            w136=> c0_n14_w136, 
            w137=> c0_n14_w137, 
            w138=> c0_n14_w138, 
            w139=> c0_n14_w139, 
            w140=> c0_n14_w140, 
            w141=> c0_n14_w141, 
            w142=> c0_n14_w142, 
            w143=> c0_n14_w143, 
            w144=> c0_n14_w144, 
            w145=> c0_n14_w145, 
            w146=> c0_n14_w146, 
            w147=> c0_n14_w147, 
            w148=> c0_n14_w148, 
            w149=> c0_n14_w149, 
            w150=> c0_n14_w150, 
            w151=> c0_n14_w151, 
            w152=> c0_n14_w152, 
            w153=> c0_n14_w153, 
            w154=> c0_n14_w154, 
            w155=> c0_n14_w155, 
            w156=> c0_n14_w156, 
            w157=> c0_n14_w157, 
            w158=> c0_n14_w158, 
            w159=> c0_n14_w159, 
            w160=> c0_n14_w160, 
            w161=> c0_n14_w161, 
            w162=> c0_n14_w162, 
            w163=> c0_n14_w163, 
            w164=> c0_n14_w164, 
            w165=> c0_n14_w165, 
            w166=> c0_n14_w166, 
            w167=> c0_n14_w167, 
            w168=> c0_n14_w168, 
            w169=> c0_n14_w169, 
            w170=> c0_n14_w170, 
            w171=> c0_n14_w171, 
            w172=> c0_n14_w172, 
            w173=> c0_n14_w173, 
            w174=> c0_n14_w174, 
            w175=> c0_n14_w175, 
            w176=> c0_n14_w176, 
            w177=> c0_n14_w177, 
            w178=> c0_n14_w178, 
            w179=> c0_n14_w179, 
            w180=> c0_n14_w180, 
            w181=> c0_n14_w181, 
            w182=> c0_n14_w182, 
            w183=> c0_n14_w183, 
            w184=> c0_n14_w184, 
            w185=> c0_n14_w185, 
            w186=> c0_n14_w186, 
            w187=> c0_n14_w187, 
            w188=> c0_n14_w188, 
            w189=> c0_n14_w189, 
            w190=> c0_n14_w190, 
            w191=> c0_n14_w191, 
            w192=> c0_n14_w192, 
            w193=> c0_n14_w193, 
            w194=> c0_n14_w194, 
            w195=> c0_n14_w195, 
            w196=> c0_n14_w196, 
            w197=> c0_n14_w197, 
            w198=> c0_n14_w198, 
            w199=> c0_n14_w199, 
            w200=> c0_n14_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n14_y
   );           
            
neuron_inst_15: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n15_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n15_w1, 
            w2=> c0_n15_w2, 
            w3=> c0_n15_w3, 
            w4=> c0_n15_w4, 
            w5=> c0_n15_w5, 
            w6=> c0_n15_w6, 
            w7=> c0_n15_w7, 
            w8=> c0_n15_w8, 
            w9=> c0_n15_w9, 
            w10=> c0_n15_w10, 
            w11=> c0_n15_w11, 
            w12=> c0_n15_w12, 
            w13=> c0_n15_w13, 
            w14=> c0_n15_w14, 
            w15=> c0_n15_w15, 
            w16=> c0_n15_w16, 
            w17=> c0_n15_w17, 
            w18=> c0_n15_w18, 
            w19=> c0_n15_w19, 
            w20=> c0_n15_w20, 
            w21=> c0_n15_w21, 
            w22=> c0_n15_w22, 
            w23=> c0_n15_w23, 
            w24=> c0_n15_w24, 
            w25=> c0_n15_w25, 
            w26=> c0_n15_w26, 
            w27=> c0_n15_w27, 
            w28=> c0_n15_w28, 
            w29=> c0_n15_w29, 
            w30=> c0_n15_w30, 
            w31=> c0_n15_w31, 
            w32=> c0_n15_w32, 
            w33=> c0_n15_w33, 
            w34=> c0_n15_w34, 
            w35=> c0_n15_w35, 
            w36=> c0_n15_w36, 
            w37=> c0_n15_w37, 
            w38=> c0_n15_w38, 
            w39=> c0_n15_w39, 
            w40=> c0_n15_w40, 
            w41=> c0_n15_w41, 
            w42=> c0_n15_w42, 
            w43=> c0_n15_w43, 
            w44=> c0_n15_w44, 
            w45=> c0_n15_w45, 
            w46=> c0_n15_w46, 
            w47=> c0_n15_w47, 
            w48=> c0_n15_w48, 
            w49=> c0_n15_w49, 
            w50=> c0_n15_w50, 
            w51=> c0_n15_w51, 
            w52=> c0_n15_w52, 
            w53=> c0_n15_w53, 
            w54=> c0_n15_w54, 
            w55=> c0_n15_w55, 
            w56=> c0_n15_w56, 
            w57=> c0_n15_w57, 
            w58=> c0_n15_w58, 
            w59=> c0_n15_w59, 
            w60=> c0_n15_w60, 
            w61=> c0_n15_w61, 
            w62=> c0_n15_w62, 
            w63=> c0_n15_w63, 
            w64=> c0_n15_w64, 
            w65=> c0_n15_w65, 
            w66=> c0_n15_w66, 
            w67=> c0_n15_w67, 
            w68=> c0_n15_w68, 
            w69=> c0_n15_w69, 
            w70=> c0_n15_w70, 
            w71=> c0_n15_w71, 
            w72=> c0_n15_w72, 
            w73=> c0_n15_w73, 
            w74=> c0_n15_w74, 
            w75=> c0_n15_w75, 
            w76=> c0_n15_w76, 
            w77=> c0_n15_w77, 
            w78=> c0_n15_w78, 
            w79=> c0_n15_w79, 
            w80=> c0_n15_w80, 
            w81=> c0_n15_w81, 
            w82=> c0_n15_w82, 
            w83=> c0_n15_w83, 
            w84=> c0_n15_w84, 
            w85=> c0_n15_w85, 
            w86=> c0_n15_w86, 
            w87=> c0_n15_w87, 
            w88=> c0_n15_w88, 
            w89=> c0_n15_w89, 
            w90=> c0_n15_w90, 
            w91=> c0_n15_w91, 
            w92=> c0_n15_w92, 
            w93=> c0_n15_w93, 
            w94=> c0_n15_w94, 
            w95=> c0_n15_w95, 
            w96=> c0_n15_w96, 
            w97=> c0_n15_w97, 
            w98=> c0_n15_w98, 
            w99=> c0_n15_w99, 
            w100=> c0_n15_w100, 
            w101=> c0_n15_w101, 
            w102=> c0_n15_w102, 
            w103=> c0_n15_w103, 
            w104=> c0_n15_w104, 
            w105=> c0_n15_w105, 
            w106=> c0_n15_w106, 
            w107=> c0_n15_w107, 
            w108=> c0_n15_w108, 
            w109=> c0_n15_w109, 
            w110=> c0_n15_w110, 
            w111=> c0_n15_w111, 
            w112=> c0_n15_w112, 
            w113=> c0_n15_w113, 
            w114=> c0_n15_w114, 
            w115=> c0_n15_w115, 
            w116=> c0_n15_w116, 
            w117=> c0_n15_w117, 
            w118=> c0_n15_w118, 
            w119=> c0_n15_w119, 
            w120=> c0_n15_w120, 
            w121=> c0_n15_w121, 
            w122=> c0_n15_w122, 
            w123=> c0_n15_w123, 
            w124=> c0_n15_w124, 
            w125=> c0_n15_w125, 
            w126=> c0_n15_w126, 
            w127=> c0_n15_w127, 
            w128=> c0_n15_w128, 
            w129=> c0_n15_w129, 
            w130=> c0_n15_w130, 
            w131=> c0_n15_w131, 
            w132=> c0_n15_w132, 
            w133=> c0_n15_w133, 
            w134=> c0_n15_w134, 
            w135=> c0_n15_w135, 
            w136=> c0_n15_w136, 
            w137=> c0_n15_w137, 
            w138=> c0_n15_w138, 
            w139=> c0_n15_w139, 
            w140=> c0_n15_w140, 
            w141=> c0_n15_w141, 
            w142=> c0_n15_w142, 
            w143=> c0_n15_w143, 
            w144=> c0_n15_w144, 
            w145=> c0_n15_w145, 
            w146=> c0_n15_w146, 
            w147=> c0_n15_w147, 
            w148=> c0_n15_w148, 
            w149=> c0_n15_w149, 
            w150=> c0_n15_w150, 
            w151=> c0_n15_w151, 
            w152=> c0_n15_w152, 
            w153=> c0_n15_w153, 
            w154=> c0_n15_w154, 
            w155=> c0_n15_w155, 
            w156=> c0_n15_w156, 
            w157=> c0_n15_w157, 
            w158=> c0_n15_w158, 
            w159=> c0_n15_w159, 
            w160=> c0_n15_w160, 
            w161=> c0_n15_w161, 
            w162=> c0_n15_w162, 
            w163=> c0_n15_w163, 
            w164=> c0_n15_w164, 
            w165=> c0_n15_w165, 
            w166=> c0_n15_w166, 
            w167=> c0_n15_w167, 
            w168=> c0_n15_w168, 
            w169=> c0_n15_w169, 
            w170=> c0_n15_w170, 
            w171=> c0_n15_w171, 
            w172=> c0_n15_w172, 
            w173=> c0_n15_w173, 
            w174=> c0_n15_w174, 
            w175=> c0_n15_w175, 
            w176=> c0_n15_w176, 
            w177=> c0_n15_w177, 
            w178=> c0_n15_w178, 
            w179=> c0_n15_w179, 
            w180=> c0_n15_w180, 
            w181=> c0_n15_w181, 
            w182=> c0_n15_w182, 
            w183=> c0_n15_w183, 
            w184=> c0_n15_w184, 
            w185=> c0_n15_w185, 
            w186=> c0_n15_w186, 
            w187=> c0_n15_w187, 
            w188=> c0_n15_w188, 
            w189=> c0_n15_w189, 
            w190=> c0_n15_w190, 
            w191=> c0_n15_w191, 
            w192=> c0_n15_w192, 
            w193=> c0_n15_w193, 
            w194=> c0_n15_w194, 
            w195=> c0_n15_w195, 
            w196=> c0_n15_w196, 
            w197=> c0_n15_w197, 
            w198=> c0_n15_w198, 
            w199=> c0_n15_w199, 
            w200=> c0_n15_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n15_y
   );           
            
neuron_inst_16: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n16_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n16_w1, 
            w2=> c0_n16_w2, 
            w3=> c0_n16_w3, 
            w4=> c0_n16_w4, 
            w5=> c0_n16_w5, 
            w6=> c0_n16_w6, 
            w7=> c0_n16_w7, 
            w8=> c0_n16_w8, 
            w9=> c0_n16_w9, 
            w10=> c0_n16_w10, 
            w11=> c0_n16_w11, 
            w12=> c0_n16_w12, 
            w13=> c0_n16_w13, 
            w14=> c0_n16_w14, 
            w15=> c0_n16_w15, 
            w16=> c0_n16_w16, 
            w17=> c0_n16_w17, 
            w18=> c0_n16_w18, 
            w19=> c0_n16_w19, 
            w20=> c0_n16_w20, 
            w21=> c0_n16_w21, 
            w22=> c0_n16_w22, 
            w23=> c0_n16_w23, 
            w24=> c0_n16_w24, 
            w25=> c0_n16_w25, 
            w26=> c0_n16_w26, 
            w27=> c0_n16_w27, 
            w28=> c0_n16_w28, 
            w29=> c0_n16_w29, 
            w30=> c0_n16_w30, 
            w31=> c0_n16_w31, 
            w32=> c0_n16_w32, 
            w33=> c0_n16_w33, 
            w34=> c0_n16_w34, 
            w35=> c0_n16_w35, 
            w36=> c0_n16_w36, 
            w37=> c0_n16_w37, 
            w38=> c0_n16_w38, 
            w39=> c0_n16_w39, 
            w40=> c0_n16_w40, 
            w41=> c0_n16_w41, 
            w42=> c0_n16_w42, 
            w43=> c0_n16_w43, 
            w44=> c0_n16_w44, 
            w45=> c0_n16_w45, 
            w46=> c0_n16_w46, 
            w47=> c0_n16_w47, 
            w48=> c0_n16_w48, 
            w49=> c0_n16_w49, 
            w50=> c0_n16_w50, 
            w51=> c0_n16_w51, 
            w52=> c0_n16_w52, 
            w53=> c0_n16_w53, 
            w54=> c0_n16_w54, 
            w55=> c0_n16_w55, 
            w56=> c0_n16_w56, 
            w57=> c0_n16_w57, 
            w58=> c0_n16_w58, 
            w59=> c0_n16_w59, 
            w60=> c0_n16_w60, 
            w61=> c0_n16_w61, 
            w62=> c0_n16_w62, 
            w63=> c0_n16_w63, 
            w64=> c0_n16_w64, 
            w65=> c0_n16_w65, 
            w66=> c0_n16_w66, 
            w67=> c0_n16_w67, 
            w68=> c0_n16_w68, 
            w69=> c0_n16_w69, 
            w70=> c0_n16_w70, 
            w71=> c0_n16_w71, 
            w72=> c0_n16_w72, 
            w73=> c0_n16_w73, 
            w74=> c0_n16_w74, 
            w75=> c0_n16_w75, 
            w76=> c0_n16_w76, 
            w77=> c0_n16_w77, 
            w78=> c0_n16_w78, 
            w79=> c0_n16_w79, 
            w80=> c0_n16_w80, 
            w81=> c0_n16_w81, 
            w82=> c0_n16_w82, 
            w83=> c0_n16_w83, 
            w84=> c0_n16_w84, 
            w85=> c0_n16_w85, 
            w86=> c0_n16_w86, 
            w87=> c0_n16_w87, 
            w88=> c0_n16_w88, 
            w89=> c0_n16_w89, 
            w90=> c0_n16_w90, 
            w91=> c0_n16_w91, 
            w92=> c0_n16_w92, 
            w93=> c0_n16_w93, 
            w94=> c0_n16_w94, 
            w95=> c0_n16_w95, 
            w96=> c0_n16_w96, 
            w97=> c0_n16_w97, 
            w98=> c0_n16_w98, 
            w99=> c0_n16_w99, 
            w100=> c0_n16_w100, 
            w101=> c0_n16_w101, 
            w102=> c0_n16_w102, 
            w103=> c0_n16_w103, 
            w104=> c0_n16_w104, 
            w105=> c0_n16_w105, 
            w106=> c0_n16_w106, 
            w107=> c0_n16_w107, 
            w108=> c0_n16_w108, 
            w109=> c0_n16_w109, 
            w110=> c0_n16_w110, 
            w111=> c0_n16_w111, 
            w112=> c0_n16_w112, 
            w113=> c0_n16_w113, 
            w114=> c0_n16_w114, 
            w115=> c0_n16_w115, 
            w116=> c0_n16_w116, 
            w117=> c0_n16_w117, 
            w118=> c0_n16_w118, 
            w119=> c0_n16_w119, 
            w120=> c0_n16_w120, 
            w121=> c0_n16_w121, 
            w122=> c0_n16_w122, 
            w123=> c0_n16_w123, 
            w124=> c0_n16_w124, 
            w125=> c0_n16_w125, 
            w126=> c0_n16_w126, 
            w127=> c0_n16_w127, 
            w128=> c0_n16_w128, 
            w129=> c0_n16_w129, 
            w130=> c0_n16_w130, 
            w131=> c0_n16_w131, 
            w132=> c0_n16_w132, 
            w133=> c0_n16_w133, 
            w134=> c0_n16_w134, 
            w135=> c0_n16_w135, 
            w136=> c0_n16_w136, 
            w137=> c0_n16_w137, 
            w138=> c0_n16_w138, 
            w139=> c0_n16_w139, 
            w140=> c0_n16_w140, 
            w141=> c0_n16_w141, 
            w142=> c0_n16_w142, 
            w143=> c0_n16_w143, 
            w144=> c0_n16_w144, 
            w145=> c0_n16_w145, 
            w146=> c0_n16_w146, 
            w147=> c0_n16_w147, 
            w148=> c0_n16_w148, 
            w149=> c0_n16_w149, 
            w150=> c0_n16_w150, 
            w151=> c0_n16_w151, 
            w152=> c0_n16_w152, 
            w153=> c0_n16_w153, 
            w154=> c0_n16_w154, 
            w155=> c0_n16_w155, 
            w156=> c0_n16_w156, 
            w157=> c0_n16_w157, 
            w158=> c0_n16_w158, 
            w159=> c0_n16_w159, 
            w160=> c0_n16_w160, 
            w161=> c0_n16_w161, 
            w162=> c0_n16_w162, 
            w163=> c0_n16_w163, 
            w164=> c0_n16_w164, 
            w165=> c0_n16_w165, 
            w166=> c0_n16_w166, 
            w167=> c0_n16_w167, 
            w168=> c0_n16_w168, 
            w169=> c0_n16_w169, 
            w170=> c0_n16_w170, 
            w171=> c0_n16_w171, 
            w172=> c0_n16_w172, 
            w173=> c0_n16_w173, 
            w174=> c0_n16_w174, 
            w175=> c0_n16_w175, 
            w176=> c0_n16_w176, 
            w177=> c0_n16_w177, 
            w178=> c0_n16_w178, 
            w179=> c0_n16_w179, 
            w180=> c0_n16_w180, 
            w181=> c0_n16_w181, 
            w182=> c0_n16_w182, 
            w183=> c0_n16_w183, 
            w184=> c0_n16_w184, 
            w185=> c0_n16_w185, 
            w186=> c0_n16_w186, 
            w187=> c0_n16_w187, 
            w188=> c0_n16_w188, 
            w189=> c0_n16_w189, 
            w190=> c0_n16_w190, 
            w191=> c0_n16_w191, 
            w192=> c0_n16_w192, 
            w193=> c0_n16_w193, 
            w194=> c0_n16_w194, 
            w195=> c0_n16_w195, 
            w196=> c0_n16_w196, 
            w197=> c0_n16_w197, 
            w198=> c0_n16_w198, 
            w199=> c0_n16_w199, 
            w200=> c0_n16_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n16_y
   );           
            
neuron_inst_17: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n17_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n17_w1, 
            w2=> c0_n17_w2, 
            w3=> c0_n17_w3, 
            w4=> c0_n17_w4, 
            w5=> c0_n17_w5, 
            w6=> c0_n17_w6, 
            w7=> c0_n17_w7, 
            w8=> c0_n17_w8, 
            w9=> c0_n17_w9, 
            w10=> c0_n17_w10, 
            w11=> c0_n17_w11, 
            w12=> c0_n17_w12, 
            w13=> c0_n17_w13, 
            w14=> c0_n17_w14, 
            w15=> c0_n17_w15, 
            w16=> c0_n17_w16, 
            w17=> c0_n17_w17, 
            w18=> c0_n17_w18, 
            w19=> c0_n17_w19, 
            w20=> c0_n17_w20, 
            w21=> c0_n17_w21, 
            w22=> c0_n17_w22, 
            w23=> c0_n17_w23, 
            w24=> c0_n17_w24, 
            w25=> c0_n17_w25, 
            w26=> c0_n17_w26, 
            w27=> c0_n17_w27, 
            w28=> c0_n17_w28, 
            w29=> c0_n17_w29, 
            w30=> c0_n17_w30, 
            w31=> c0_n17_w31, 
            w32=> c0_n17_w32, 
            w33=> c0_n17_w33, 
            w34=> c0_n17_w34, 
            w35=> c0_n17_w35, 
            w36=> c0_n17_w36, 
            w37=> c0_n17_w37, 
            w38=> c0_n17_w38, 
            w39=> c0_n17_w39, 
            w40=> c0_n17_w40, 
            w41=> c0_n17_w41, 
            w42=> c0_n17_w42, 
            w43=> c0_n17_w43, 
            w44=> c0_n17_w44, 
            w45=> c0_n17_w45, 
            w46=> c0_n17_w46, 
            w47=> c0_n17_w47, 
            w48=> c0_n17_w48, 
            w49=> c0_n17_w49, 
            w50=> c0_n17_w50, 
            w51=> c0_n17_w51, 
            w52=> c0_n17_w52, 
            w53=> c0_n17_w53, 
            w54=> c0_n17_w54, 
            w55=> c0_n17_w55, 
            w56=> c0_n17_w56, 
            w57=> c0_n17_w57, 
            w58=> c0_n17_w58, 
            w59=> c0_n17_w59, 
            w60=> c0_n17_w60, 
            w61=> c0_n17_w61, 
            w62=> c0_n17_w62, 
            w63=> c0_n17_w63, 
            w64=> c0_n17_w64, 
            w65=> c0_n17_w65, 
            w66=> c0_n17_w66, 
            w67=> c0_n17_w67, 
            w68=> c0_n17_w68, 
            w69=> c0_n17_w69, 
            w70=> c0_n17_w70, 
            w71=> c0_n17_w71, 
            w72=> c0_n17_w72, 
            w73=> c0_n17_w73, 
            w74=> c0_n17_w74, 
            w75=> c0_n17_w75, 
            w76=> c0_n17_w76, 
            w77=> c0_n17_w77, 
            w78=> c0_n17_w78, 
            w79=> c0_n17_w79, 
            w80=> c0_n17_w80, 
            w81=> c0_n17_w81, 
            w82=> c0_n17_w82, 
            w83=> c0_n17_w83, 
            w84=> c0_n17_w84, 
            w85=> c0_n17_w85, 
            w86=> c0_n17_w86, 
            w87=> c0_n17_w87, 
            w88=> c0_n17_w88, 
            w89=> c0_n17_w89, 
            w90=> c0_n17_w90, 
            w91=> c0_n17_w91, 
            w92=> c0_n17_w92, 
            w93=> c0_n17_w93, 
            w94=> c0_n17_w94, 
            w95=> c0_n17_w95, 
            w96=> c0_n17_w96, 
            w97=> c0_n17_w97, 
            w98=> c0_n17_w98, 
            w99=> c0_n17_w99, 
            w100=> c0_n17_w100, 
            w101=> c0_n17_w101, 
            w102=> c0_n17_w102, 
            w103=> c0_n17_w103, 
            w104=> c0_n17_w104, 
            w105=> c0_n17_w105, 
            w106=> c0_n17_w106, 
            w107=> c0_n17_w107, 
            w108=> c0_n17_w108, 
            w109=> c0_n17_w109, 
            w110=> c0_n17_w110, 
            w111=> c0_n17_w111, 
            w112=> c0_n17_w112, 
            w113=> c0_n17_w113, 
            w114=> c0_n17_w114, 
            w115=> c0_n17_w115, 
            w116=> c0_n17_w116, 
            w117=> c0_n17_w117, 
            w118=> c0_n17_w118, 
            w119=> c0_n17_w119, 
            w120=> c0_n17_w120, 
            w121=> c0_n17_w121, 
            w122=> c0_n17_w122, 
            w123=> c0_n17_w123, 
            w124=> c0_n17_w124, 
            w125=> c0_n17_w125, 
            w126=> c0_n17_w126, 
            w127=> c0_n17_w127, 
            w128=> c0_n17_w128, 
            w129=> c0_n17_w129, 
            w130=> c0_n17_w130, 
            w131=> c0_n17_w131, 
            w132=> c0_n17_w132, 
            w133=> c0_n17_w133, 
            w134=> c0_n17_w134, 
            w135=> c0_n17_w135, 
            w136=> c0_n17_w136, 
            w137=> c0_n17_w137, 
            w138=> c0_n17_w138, 
            w139=> c0_n17_w139, 
            w140=> c0_n17_w140, 
            w141=> c0_n17_w141, 
            w142=> c0_n17_w142, 
            w143=> c0_n17_w143, 
            w144=> c0_n17_w144, 
            w145=> c0_n17_w145, 
            w146=> c0_n17_w146, 
            w147=> c0_n17_w147, 
            w148=> c0_n17_w148, 
            w149=> c0_n17_w149, 
            w150=> c0_n17_w150, 
            w151=> c0_n17_w151, 
            w152=> c0_n17_w152, 
            w153=> c0_n17_w153, 
            w154=> c0_n17_w154, 
            w155=> c0_n17_w155, 
            w156=> c0_n17_w156, 
            w157=> c0_n17_w157, 
            w158=> c0_n17_w158, 
            w159=> c0_n17_w159, 
            w160=> c0_n17_w160, 
            w161=> c0_n17_w161, 
            w162=> c0_n17_w162, 
            w163=> c0_n17_w163, 
            w164=> c0_n17_w164, 
            w165=> c0_n17_w165, 
            w166=> c0_n17_w166, 
            w167=> c0_n17_w167, 
            w168=> c0_n17_w168, 
            w169=> c0_n17_w169, 
            w170=> c0_n17_w170, 
            w171=> c0_n17_w171, 
            w172=> c0_n17_w172, 
            w173=> c0_n17_w173, 
            w174=> c0_n17_w174, 
            w175=> c0_n17_w175, 
            w176=> c0_n17_w176, 
            w177=> c0_n17_w177, 
            w178=> c0_n17_w178, 
            w179=> c0_n17_w179, 
            w180=> c0_n17_w180, 
            w181=> c0_n17_w181, 
            w182=> c0_n17_w182, 
            w183=> c0_n17_w183, 
            w184=> c0_n17_w184, 
            w185=> c0_n17_w185, 
            w186=> c0_n17_w186, 
            w187=> c0_n17_w187, 
            w188=> c0_n17_w188, 
            w189=> c0_n17_w189, 
            w190=> c0_n17_w190, 
            w191=> c0_n17_w191, 
            w192=> c0_n17_w192, 
            w193=> c0_n17_w193, 
            w194=> c0_n17_w194, 
            w195=> c0_n17_w195, 
            w196=> c0_n17_w196, 
            w197=> c0_n17_w197, 
            w198=> c0_n17_w198, 
            w199=> c0_n17_w199, 
            w200=> c0_n17_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n17_y
   );           
            
neuron_inst_18: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n18_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n18_w1, 
            w2=> c0_n18_w2, 
            w3=> c0_n18_w3, 
            w4=> c0_n18_w4, 
            w5=> c0_n18_w5, 
            w6=> c0_n18_w6, 
            w7=> c0_n18_w7, 
            w8=> c0_n18_w8, 
            w9=> c0_n18_w9, 
            w10=> c0_n18_w10, 
            w11=> c0_n18_w11, 
            w12=> c0_n18_w12, 
            w13=> c0_n18_w13, 
            w14=> c0_n18_w14, 
            w15=> c0_n18_w15, 
            w16=> c0_n18_w16, 
            w17=> c0_n18_w17, 
            w18=> c0_n18_w18, 
            w19=> c0_n18_w19, 
            w20=> c0_n18_w20, 
            w21=> c0_n18_w21, 
            w22=> c0_n18_w22, 
            w23=> c0_n18_w23, 
            w24=> c0_n18_w24, 
            w25=> c0_n18_w25, 
            w26=> c0_n18_w26, 
            w27=> c0_n18_w27, 
            w28=> c0_n18_w28, 
            w29=> c0_n18_w29, 
            w30=> c0_n18_w30, 
            w31=> c0_n18_w31, 
            w32=> c0_n18_w32, 
            w33=> c0_n18_w33, 
            w34=> c0_n18_w34, 
            w35=> c0_n18_w35, 
            w36=> c0_n18_w36, 
            w37=> c0_n18_w37, 
            w38=> c0_n18_w38, 
            w39=> c0_n18_w39, 
            w40=> c0_n18_w40, 
            w41=> c0_n18_w41, 
            w42=> c0_n18_w42, 
            w43=> c0_n18_w43, 
            w44=> c0_n18_w44, 
            w45=> c0_n18_w45, 
            w46=> c0_n18_w46, 
            w47=> c0_n18_w47, 
            w48=> c0_n18_w48, 
            w49=> c0_n18_w49, 
            w50=> c0_n18_w50, 
            w51=> c0_n18_w51, 
            w52=> c0_n18_w52, 
            w53=> c0_n18_w53, 
            w54=> c0_n18_w54, 
            w55=> c0_n18_w55, 
            w56=> c0_n18_w56, 
            w57=> c0_n18_w57, 
            w58=> c0_n18_w58, 
            w59=> c0_n18_w59, 
            w60=> c0_n18_w60, 
            w61=> c0_n18_w61, 
            w62=> c0_n18_w62, 
            w63=> c0_n18_w63, 
            w64=> c0_n18_w64, 
            w65=> c0_n18_w65, 
            w66=> c0_n18_w66, 
            w67=> c0_n18_w67, 
            w68=> c0_n18_w68, 
            w69=> c0_n18_w69, 
            w70=> c0_n18_w70, 
            w71=> c0_n18_w71, 
            w72=> c0_n18_w72, 
            w73=> c0_n18_w73, 
            w74=> c0_n18_w74, 
            w75=> c0_n18_w75, 
            w76=> c0_n18_w76, 
            w77=> c0_n18_w77, 
            w78=> c0_n18_w78, 
            w79=> c0_n18_w79, 
            w80=> c0_n18_w80, 
            w81=> c0_n18_w81, 
            w82=> c0_n18_w82, 
            w83=> c0_n18_w83, 
            w84=> c0_n18_w84, 
            w85=> c0_n18_w85, 
            w86=> c0_n18_w86, 
            w87=> c0_n18_w87, 
            w88=> c0_n18_w88, 
            w89=> c0_n18_w89, 
            w90=> c0_n18_w90, 
            w91=> c0_n18_w91, 
            w92=> c0_n18_w92, 
            w93=> c0_n18_w93, 
            w94=> c0_n18_w94, 
            w95=> c0_n18_w95, 
            w96=> c0_n18_w96, 
            w97=> c0_n18_w97, 
            w98=> c0_n18_w98, 
            w99=> c0_n18_w99, 
            w100=> c0_n18_w100, 
            w101=> c0_n18_w101, 
            w102=> c0_n18_w102, 
            w103=> c0_n18_w103, 
            w104=> c0_n18_w104, 
            w105=> c0_n18_w105, 
            w106=> c0_n18_w106, 
            w107=> c0_n18_w107, 
            w108=> c0_n18_w108, 
            w109=> c0_n18_w109, 
            w110=> c0_n18_w110, 
            w111=> c0_n18_w111, 
            w112=> c0_n18_w112, 
            w113=> c0_n18_w113, 
            w114=> c0_n18_w114, 
            w115=> c0_n18_w115, 
            w116=> c0_n18_w116, 
            w117=> c0_n18_w117, 
            w118=> c0_n18_w118, 
            w119=> c0_n18_w119, 
            w120=> c0_n18_w120, 
            w121=> c0_n18_w121, 
            w122=> c0_n18_w122, 
            w123=> c0_n18_w123, 
            w124=> c0_n18_w124, 
            w125=> c0_n18_w125, 
            w126=> c0_n18_w126, 
            w127=> c0_n18_w127, 
            w128=> c0_n18_w128, 
            w129=> c0_n18_w129, 
            w130=> c0_n18_w130, 
            w131=> c0_n18_w131, 
            w132=> c0_n18_w132, 
            w133=> c0_n18_w133, 
            w134=> c0_n18_w134, 
            w135=> c0_n18_w135, 
            w136=> c0_n18_w136, 
            w137=> c0_n18_w137, 
            w138=> c0_n18_w138, 
            w139=> c0_n18_w139, 
            w140=> c0_n18_w140, 
            w141=> c0_n18_w141, 
            w142=> c0_n18_w142, 
            w143=> c0_n18_w143, 
            w144=> c0_n18_w144, 
            w145=> c0_n18_w145, 
            w146=> c0_n18_w146, 
            w147=> c0_n18_w147, 
            w148=> c0_n18_w148, 
            w149=> c0_n18_w149, 
            w150=> c0_n18_w150, 
            w151=> c0_n18_w151, 
            w152=> c0_n18_w152, 
            w153=> c0_n18_w153, 
            w154=> c0_n18_w154, 
            w155=> c0_n18_w155, 
            w156=> c0_n18_w156, 
            w157=> c0_n18_w157, 
            w158=> c0_n18_w158, 
            w159=> c0_n18_w159, 
            w160=> c0_n18_w160, 
            w161=> c0_n18_w161, 
            w162=> c0_n18_w162, 
            w163=> c0_n18_w163, 
            w164=> c0_n18_w164, 
            w165=> c0_n18_w165, 
            w166=> c0_n18_w166, 
            w167=> c0_n18_w167, 
            w168=> c0_n18_w168, 
            w169=> c0_n18_w169, 
            w170=> c0_n18_w170, 
            w171=> c0_n18_w171, 
            w172=> c0_n18_w172, 
            w173=> c0_n18_w173, 
            w174=> c0_n18_w174, 
            w175=> c0_n18_w175, 
            w176=> c0_n18_w176, 
            w177=> c0_n18_w177, 
            w178=> c0_n18_w178, 
            w179=> c0_n18_w179, 
            w180=> c0_n18_w180, 
            w181=> c0_n18_w181, 
            w182=> c0_n18_w182, 
            w183=> c0_n18_w183, 
            w184=> c0_n18_w184, 
            w185=> c0_n18_w185, 
            w186=> c0_n18_w186, 
            w187=> c0_n18_w187, 
            w188=> c0_n18_w188, 
            w189=> c0_n18_w189, 
            w190=> c0_n18_w190, 
            w191=> c0_n18_w191, 
            w192=> c0_n18_w192, 
            w193=> c0_n18_w193, 
            w194=> c0_n18_w194, 
            w195=> c0_n18_w195, 
            w196=> c0_n18_w196, 
            w197=> c0_n18_w197, 
            w198=> c0_n18_w198, 
            w199=> c0_n18_w199, 
            w200=> c0_n18_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n18_y
   );           
            
neuron_inst_19: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n19_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n19_w1, 
            w2=> c0_n19_w2, 
            w3=> c0_n19_w3, 
            w4=> c0_n19_w4, 
            w5=> c0_n19_w5, 
            w6=> c0_n19_w6, 
            w7=> c0_n19_w7, 
            w8=> c0_n19_w8, 
            w9=> c0_n19_w9, 
            w10=> c0_n19_w10, 
            w11=> c0_n19_w11, 
            w12=> c0_n19_w12, 
            w13=> c0_n19_w13, 
            w14=> c0_n19_w14, 
            w15=> c0_n19_w15, 
            w16=> c0_n19_w16, 
            w17=> c0_n19_w17, 
            w18=> c0_n19_w18, 
            w19=> c0_n19_w19, 
            w20=> c0_n19_w20, 
            w21=> c0_n19_w21, 
            w22=> c0_n19_w22, 
            w23=> c0_n19_w23, 
            w24=> c0_n19_w24, 
            w25=> c0_n19_w25, 
            w26=> c0_n19_w26, 
            w27=> c0_n19_w27, 
            w28=> c0_n19_w28, 
            w29=> c0_n19_w29, 
            w30=> c0_n19_w30, 
            w31=> c0_n19_w31, 
            w32=> c0_n19_w32, 
            w33=> c0_n19_w33, 
            w34=> c0_n19_w34, 
            w35=> c0_n19_w35, 
            w36=> c0_n19_w36, 
            w37=> c0_n19_w37, 
            w38=> c0_n19_w38, 
            w39=> c0_n19_w39, 
            w40=> c0_n19_w40, 
            w41=> c0_n19_w41, 
            w42=> c0_n19_w42, 
            w43=> c0_n19_w43, 
            w44=> c0_n19_w44, 
            w45=> c0_n19_w45, 
            w46=> c0_n19_w46, 
            w47=> c0_n19_w47, 
            w48=> c0_n19_w48, 
            w49=> c0_n19_w49, 
            w50=> c0_n19_w50, 
            w51=> c0_n19_w51, 
            w52=> c0_n19_w52, 
            w53=> c0_n19_w53, 
            w54=> c0_n19_w54, 
            w55=> c0_n19_w55, 
            w56=> c0_n19_w56, 
            w57=> c0_n19_w57, 
            w58=> c0_n19_w58, 
            w59=> c0_n19_w59, 
            w60=> c0_n19_w60, 
            w61=> c0_n19_w61, 
            w62=> c0_n19_w62, 
            w63=> c0_n19_w63, 
            w64=> c0_n19_w64, 
            w65=> c0_n19_w65, 
            w66=> c0_n19_w66, 
            w67=> c0_n19_w67, 
            w68=> c0_n19_w68, 
            w69=> c0_n19_w69, 
            w70=> c0_n19_w70, 
            w71=> c0_n19_w71, 
            w72=> c0_n19_w72, 
            w73=> c0_n19_w73, 
            w74=> c0_n19_w74, 
            w75=> c0_n19_w75, 
            w76=> c0_n19_w76, 
            w77=> c0_n19_w77, 
            w78=> c0_n19_w78, 
            w79=> c0_n19_w79, 
            w80=> c0_n19_w80, 
            w81=> c0_n19_w81, 
            w82=> c0_n19_w82, 
            w83=> c0_n19_w83, 
            w84=> c0_n19_w84, 
            w85=> c0_n19_w85, 
            w86=> c0_n19_w86, 
            w87=> c0_n19_w87, 
            w88=> c0_n19_w88, 
            w89=> c0_n19_w89, 
            w90=> c0_n19_w90, 
            w91=> c0_n19_w91, 
            w92=> c0_n19_w92, 
            w93=> c0_n19_w93, 
            w94=> c0_n19_w94, 
            w95=> c0_n19_w95, 
            w96=> c0_n19_w96, 
            w97=> c0_n19_w97, 
            w98=> c0_n19_w98, 
            w99=> c0_n19_w99, 
            w100=> c0_n19_w100, 
            w101=> c0_n19_w101, 
            w102=> c0_n19_w102, 
            w103=> c0_n19_w103, 
            w104=> c0_n19_w104, 
            w105=> c0_n19_w105, 
            w106=> c0_n19_w106, 
            w107=> c0_n19_w107, 
            w108=> c0_n19_w108, 
            w109=> c0_n19_w109, 
            w110=> c0_n19_w110, 
            w111=> c0_n19_w111, 
            w112=> c0_n19_w112, 
            w113=> c0_n19_w113, 
            w114=> c0_n19_w114, 
            w115=> c0_n19_w115, 
            w116=> c0_n19_w116, 
            w117=> c0_n19_w117, 
            w118=> c0_n19_w118, 
            w119=> c0_n19_w119, 
            w120=> c0_n19_w120, 
            w121=> c0_n19_w121, 
            w122=> c0_n19_w122, 
            w123=> c0_n19_w123, 
            w124=> c0_n19_w124, 
            w125=> c0_n19_w125, 
            w126=> c0_n19_w126, 
            w127=> c0_n19_w127, 
            w128=> c0_n19_w128, 
            w129=> c0_n19_w129, 
            w130=> c0_n19_w130, 
            w131=> c0_n19_w131, 
            w132=> c0_n19_w132, 
            w133=> c0_n19_w133, 
            w134=> c0_n19_w134, 
            w135=> c0_n19_w135, 
            w136=> c0_n19_w136, 
            w137=> c0_n19_w137, 
            w138=> c0_n19_w138, 
            w139=> c0_n19_w139, 
            w140=> c0_n19_w140, 
            w141=> c0_n19_w141, 
            w142=> c0_n19_w142, 
            w143=> c0_n19_w143, 
            w144=> c0_n19_w144, 
            w145=> c0_n19_w145, 
            w146=> c0_n19_w146, 
            w147=> c0_n19_w147, 
            w148=> c0_n19_w148, 
            w149=> c0_n19_w149, 
            w150=> c0_n19_w150, 
            w151=> c0_n19_w151, 
            w152=> c0_n19_w152, 
            w153=> c0_n19_w153, 
            w154=> c0_n19_w154, 
            w155=> c0_n19_w155, 
            w156=> c0_n19_w156, 
            w157=> c0_n19_w157, 
            w158=> c0_n19_w158, 
            w159=> c0_n19_w159, 
            w160=> c0_n19_w160, 
            w161=> c0_n19_w161, 
            w162=> c0_n19_w162, 
            w163=> c0_n19_w163, 
            w164=> c0_n19_w164, 
            w165=> c0_n19_w165, 
            w166=> c0_n19_w166, 
            w167=> c0_n19_w167, 
            w168=> c0_n19_w168, 
            w169=> c0_n19_w169, 
            w170=> c0_n19_w170, 
            w171=> c0_n19_w171, 
            w172=> c0_n19_w172, 
            w173=> c0_n19_w173, 
            w174=> c0_n19_w174, 
            w175=> c0_n19_w175, 
            w176=> c0_n19_w176, 
            w177=> c0_n19_w177, 
            w178=> c0_n19_w178, 
            w179=> c0_n19_w179, 
            w180=> c0_n19_w180, 
            w181=> c0_n19_w181, 
            w182=> c0_n19_w182, 
            w183=> c0_n19_w183, 
            w184=> c0_n19_w184, 
            w185=> c0_n19_w185, 
            w186=> c0_n19_w186, 
            w187=> c0_n19_w187, 
            w188=> c0_n19_w188, 
            w189=> c0_n19_w189, 
            w190=> c0_n19_w190, 
            w191=> c0_n19_w191, 
            w192=> c0_n19_w192, 
            w193=> c0_n19_w193, 
            w194=> c0_n19_w194, 
            w195=> c0_n19_w195, 
            w196=> c0_n19_w196, 
            w197=> c0_n19_w197, 
            w198=> c0_n19_w198, 
            w199=> c0_n19_w199, 
            w200=> c0_n19_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n19_y
   );           
            
neuron_inst_20: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n20_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n20_w1, 
            w2=> c0_n20_w2, 
            w3=> c0_n20_w3, 
            w4=> c0_n20_w4, 
            w5=> c0_n20_w5, 
            w6=> c0_n20_w6, 
            w7=> c0_n20_w7, 
            w8=> c0_n20_w8, 
            w9=> c0_n20_w9, 
            w10=> c0_n20_w10, 
            w11=> c0_n20_w11, 
            w12=> c0_n20_w12, 
            w13=> c0_n20_w13, 
            w14=> c0_n20_w14, 
            w15=> c0_n20_w15, 
            w16=> c0_n20_w16, 
            w17=> c0_n20_w17, 
            w18=> c0_n20_w18, 
            w19=> c0_n20_w19, 
            w20=> c0_n20_w20, 
            w21=> c0_n20_w21, 
            w22=> c0_n20_w22, 
            w23=> c0_n20_w23, 
            w24=> c0_n20_w24, 
            w25=> c0_n20_w25, 
            w26=> c0_n20_w26, 
            w27=> c0_n20_w27, 
            w28=> c0_n20_w28, 
            w29=> c0_n20_w29, 
            w30=> c0_n20_w30, 
            w31=> c0_n20_w31, 
            w32=> c0_n20_w32, 
            w33=> c0_n20_w33, 
            w34=> c0_n20_w34, 
            w35=> c0_n20_w35, 
            w36=> c0_n20_w36, 
            w37=> c0_n20_w37, 
            w38=> c0_n20_w38, 
            w39=> c0_n20_w39, 
            w40=> c0_n20_w40, 
            w41=> c0_n20_w41, 
            w42=> c0_n20_w42, 
            w43=> c0_n20_w43, 
            w44=> c0_n20_w44, 
            w45=> c0_n20_w45, 
            w46=> c0_n20_w46, 
            w47=> c0_n20_w47, 
            w48=> c0_n20_w48, 
            w49=> c0_n20_w49, 
            w50=> c0_n20_w50, 
            w51=> c0_n20_w51, 
            w52=> c0_n20_w52, 
            w53=> c0_n20_w53, 
            w54=> c0_n20_w54, 
            w55=> c0_n20_w55, 
            w56=> c0_n20_w56, 
            w57=> c0_n20_w57, 
            w58=> c0_n20_w58, 
            w59=> c0_n20_w59, 
            w60=> c0_n20_w60, 
            w61=> c0_n20_w61, 
            w62=> c0_n20_w62, 
            w63=> c0_n20_w63, 
            w64=> c0_n20_w64, 
            w65=> c0_n20_w65, 
            w66=> c0_n20_w66, 
            w67=> c0_n20_w67, 
            w68=> c0_n20_w68, 
            w69=> c0_n20_w69, 
            w70=> c0_n20_w70, 
            w71=> c0_n20_w71, 
            w72=> c0_n20_w72, 
            w73=> c0_n20_w73, 
            w74=> c0_n20_w74, 
            w75=> c0_n20_w75, 
            w76=> c0_n20_w76, 
            w77=> c0_n20_w77, 
            w78=> c0_n20_w78, 
            w79=> c0_n20_w79, 
            w80=> c0_n20_w80, 
            w81=> c0_n20_w81, 
            w82=> c0_n20_w82, 
            w83=> c0_n20_w83, 
            w84=> c0_n20_w84, 
            w85=> c0_n20_w85, 
            w86=> c0_n20_w86, 
            w87=> c0_n20_w87, 
            w88=> c0_n20_w88, 
            w89=> c0_n20_w89, 
            w90=> c0_n20_w90, 
            w91=> c0_n20_w91, 
            w92=> c0_n20_w92, 
            w93=> c0_n20_w93, 
            w94=> c0_n20_w94, 
            w95=> c0_n20_w95, 
            w96=> c0_n20_w96, 
            w97=> c0_n20_w97, 
            w98=> c0_n20_w98, 
            w99=> c0_n20_w99, 
            w100=> c0_n20_w100, 
            w101=> c0_n20_w101, 
            w102=> c0_n20_w102, 
            w103=> c0_n20_w103, 
            w104=> c0_n20_w104, 
            w105=> c0_n20_w105, 
            w106=> c0_n20_w106, 
            w107=> c0_n20_w107, 
            w108=> c0_n20_w108, 
            w109=> c0_n20_w109, 
            w110=> c0_n20_w110, 
            w111=> c0_n20_w111, 
            w112=> c0_n20_w112, 
            w113=> c0_n20_w113, 
            w114=> c0_n20_w114, 
            w115=> c0_n20_w115, 
            w116=> c0_n20_w116, 
            w117=> c0_n20_w117, 
            w118=> c0_n20_w118, 
            w119=> c0_n20_w119, 
            w120=> c0_n20_w120, 
            w121=> c0_n20_w121, 
            w122=> c0_n20_w122, 
            w123=> c0_n20_w123, 
            w124=> c0_n20_w124, 
            w125=> c0_n20_w125, 
            w126=> c0_n20_w126, 
            w127=> c0_n20_w127, 
            w128=> c0_n20_w128, 
            w129=> c0_n20_w129, 
            w130=> c0_n20_w130, 
            w131=> c0_n20_w131, 
            w132=> c0_n20_w132, 
            w133=> c0_n20_w133, 
            w134=> c0_n20_w134, 
            w135=> c0_n20_w135, 
            w136=> c0_n20_w136, 
            w137=> c0_n20_w137, 
            w138=> c0_n20_w138, 
            w139=> c0_n20_w139, 
            w140=> c0_n20_w140, 
            w141=> c0_n20_w141, 
            w142=> c0_n20_w142, 
            w143=> c0_n20_w143, 
            w144=> c0_n20_w144, 
            w145=> c0_n20_w145, 
            w146=> c0_n20_w146, 
            w147=> c0_n20_w147, 
            w148=> c0_n20_w148, 
            w149=> c0_n20_w149, 
            w150=> c0_n20_w150, 
            w151=> c0_n20_w151, 
            w152=> c0_n20_w152, 
            w153=> c0_n20_w153, 
            w154=> c0_n20_w154, 
            w155=> c0_n20_w155, 
            w156=> c0_n20_w156, 
            w157=> c0_n20_w157, 
            w158=> c0_n20_w158, 
            w159=> c0_n20_w159, 
            w160=> c0_n20_w160, 
            w161=> c0_n20_w161, 
            w162=> c0_n20_w162, 
            w163=> c0_n20_w163, 
            w164=> c0_n20_w164, 
            w165=> c0_n20_w165, 
            w166=> c0_n20_w166, 
            w167=> c0_n20_w167, 
            w168=> c0_n20_w168, 
            w169=> c0_n20_w169, 
            w170=> c0_n20_w170, 
            w171=> c0_n20_w171, 
            w172=> c0_n20_w172, 
            w173=> c0_n20_w173, 
            w174=> c0_n20_w174, 
            w175=> c0_n20_w175, 
            w176=> c0_n20_w176, 
            w177=> c0_n20_w177, 
            w178=> c0_n20_w178, 
            w179=> c0_n20_w179, 
            w180=> c0_n20_w180, 
            w181=> c0_n20_w181, 
            w182=> c0_n20_w182, 
            w183=> c0_n20_w183, 
            w184=> c0_n20_w184, 
            w185=> c0_n20_w185, 
            w186=> c0_n20_w186, 
            w187=> c0_n20_w187, 
            w188=> c0_n20_w188, 
            w189=> c0_n20_w189, 
            w190=> c0_n20_w190, 
            w191=> c0_n20_w191, 
            w192=> c0_n20_w192, 
            w193=> c0_n20_w193, 
            w194=> c0_n20_w194, 
            w195=> c0_n20_w195, 
            w196=> c0_n20_w196, 
            w197=> c0_n20_w197, 
            w198=> c0_n20_w198, 
            w199=> c0_n20_w199, 
            w200=> c0_n20_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n20_y
   );           
            
neuron_inst_21: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n21_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n21_w1, 
            w2=> c0_n21_w2, 
            w3=> c0_n21_w3, 
            w4=> c0_n21_w4, 
            w5=> c0_n21_w5, 
            w6=> c0_n21_w6, 
            w7=> c0_n21_w7, 
            w8=> c0_n21_w8, 
            w9=> c0_n21_w9, 
            w10=> c0_n21_w10, 
            w11=> c0_n21_w11, 
            w12=> c0_n21_w12, 
            w13=> c0_n21_w13, 
            w14=> c0_n21_w14, 
            w15=> c0_n21_w15, 
            w16=> c0_n21_w16, 
            w17=> c0_n21_w17, 
            w18=> c0_n21_w18, 
            w19=> c0_n21_w19, 
            w20=> c0_n21_w20, 
            w21=> c0_n21_w21, 
            w22=> c0_n21_w22, 
            w23=> c0_n21_w23, 
            w24=> c0_n21_w24, 
            w25=> c0_n21_w25, 
            w26=> c0_n21_w26, 
            w27=> c0_n21_w27, 
            w28=> c0_n21_w28, 
            w29=> c0_n21_w29, 
            w30=> c0_n21_w30, 
            w31=> c0_n21_w31, 
            w32=> c0_n21_w32, 
            w33=> c0_n21_w33, 
            w34=> c0_n21_w34, 
            w35=> c0_n21_w35, 
            w36=> c0_n21_w36, 
            w37=> c0_n21_w37, 
            w38=> c0_n21_w38, 
            w39=> c0_n21_w39, 
            w40=> c0_n21_w40, 
            w41=> c0_n21_w41, 
            w42=> c0_n21_w42, 
            w43=> c0_n21_w43, 
            w44=> c0_n21_w44, 
            w45=> c0_n21_w45, 
            w46=> c0_n21_w46, 
            w47=> c0_n21_w47, 
            w48=> c0_n21_w48, 
            w49=> c0_n21_w49, 
            w50=> c0_n21_w50, 
            w51=> c0_n21_w51, 
            w52=> c0_n21_w52, 
            w53=> c0_n21_w53, 
            w54=> c0_n21_w54, 
            w55=> c0_n21_w55, 
            w56=> c0_n21_w56, 
            w57=> c0_n21_w57, 
            w58=> c0_n21_w58, 
            w59=> c0_n21_w59, 
            w60=> c0_n21_w60, 
            w61=> c0_n21_w61, 
            w62=> c0_n21_w62, 
            w63=> c0_n21_w63, 
            w64=> c0_n21_w64, 
            w65=> c0_n21_w65, 
            w66=> c0_n21_w66, 
            w67=> c0_n21_w67, 
            w68=> c0_n21_w68, 
            w69=> c0_n21_w69, 
            w70=> c0_n21_w70, 
            w71=> c0_n21_w71, 
            w72=> c0_n21_w72, 
            w73=> c0_n21_w73, 
            w74=> c0_n21_w74, 
            w75=> c0_n21_w75, 
            w76=> c0_n21_w76, 
            w77=> c0_n21_w77, 
            w78=> c0_n21_w78, 
            w79=> c0_n21_w79, 
            w80=> c0_n21_w80, 
            w81=> c0_n21_w81, 
            w82=> c0_n21_w82, 
            w83=> c0_n21_w83, 
            w84=> c0_n21_w84, 
            w85=> c0_n21_w85, 
            w86=> c0_n21_w86, 
            w87=> c0_n21_w87, 
            w88=> c0_n21_w88, 
            w89=> c0_n21_w89, 
            w90=> c0_n21_w90, 
            w91=> c0_n21_w91, 
            w92=> c0_n21_w92, 
            w93=> c0_n21_w93, 
            w94=> c0_n21_w94, 
            w95=> c0_n21_w95, 
            w96=> c0_n21_w96, 
            w97=> c0_n21_w97, 
            w98=> c0_n21_w98, 
            w99=> c0_n21_w99, 
            w100=> c0_n21_w100, 
            w101=> c0_n21_w101, 
            w102=> c0_n21_w102, 
            w103=> c0_n21_w103, 
            w104=> c0_n21_w104, 
            w105=> c0_n21_w105, 
            w106=> c0_n21_w106, 
            w107=> c0_n21_w107, 
            w108=> c0_n21_w108, 
            w109=> c0_n21_w109, 
            w110=> c0_n21_w110, 
            w111=> c0_n21_w111, 
            w112=> c0_n21_w112, 
            w113=> c0_n21_w113, 
            w114=> c0_n21_w114, 
            w115=> c0_n21_w115, 
            w116=> c0_n21_w116, 
            w117=> c0_n21_w117, 
            w118=> c0_n21_w118, 
            w119=> c0_n21_w119, 
            w120=> c0_n21_w120, 
            w121=> c0_n21_w121, 
            w122=> c0_n21_w122, 
            w123=> c0_n21_w123, 
            w124=> c0_n21_w124, 
            w125=> c0_n21_w125, 
            w126=> c0_n21_w126, 
            w127=> c0_n21_w127, 
            w128=> c0_n21_w128, 
            w129=> c0_n21_w129, 
            w130=> c0_n21_w130, 
            w131=> c0_n21_w131, 
            w132=> c0_n21_w132, 
            w133=> c0_n21_w133, 
            w134=> c0_n21_w134, 
            w135=> c0_n21_w135, 
            w136=> c0_n21_w136, 
            w137=> c0_n21_w137, 
            w138=> c0_n21_w138, 
            w139=> c0_n21_w139, 
            w140=> c0_n21_w140, 
            w141=> c0_n21_w141, 
            w142=> c0_n21_w142, 
            w143=> c0_n21_w143, 
            w144=> c0_n21_w144, 
            w145=> c0_n21_w145, 
            w146=> c0_n21_w146, 
            w147=> c0_n21_w147, 
            w148=> c0_n21_w148, 
            w149=> c0_n21_w149, 
            w150=> c0_n21_w150, 
            w151=> c0_n21_w151, 
            w152=> c0_n21_w152, 
            w153=> c0_n21_w153, 
            w154=> c0_n21_w154, 
            w155=> c0_n21_w155, 
            w156=> c0_n21_w156, 
            w157=> c0_n21_w157, 
            w158=> c0_n21_w158, 
            w159=> c0_n21_w159, 
            w160=> c0_n21_w160, 
            w161=> c0_n21_w161, 
            w162=> c0_n21_w162, 
            w163=> c0_n21_w163, 
            w164=> c0_n21_w164, 
            w165=> c0_n21_w165, 
            w166=> c0_n21_w166, 
            w167=> c0_n21_w167, 
            w168=> c0_n21_w168, 
            w169=> c0_n21_w169, 
            w170=> c0_n21_w170, 
            w171=> c0_n21_w171, 
            w172=> c0_n21_w172, 
            w173=> c0_n21_w173, 
            w174=> c0_n21_w174, 
            w175=> c0_n21_w175, 
            w176=> c0_n21_w176, 
            w177=> c0_n21_w177, 
            w178=> c0_n21_w178, 
            w179=> c0_n21_w179, 
            w180=> c0_n21_w180, 
            w181=> c0_n21_w181, 
            w182=> c0_n21_w182, 
            w183=> c0_n21_w183, 
            w184=> c0_n21_w184, 
            w185=> c0_n21_w185, 
            w186=> c0_n21_w186, 
            w187=> c0_n21_w187, 
            w188=> c0_n21_w188, 
            w189=> c0_n21_w189, 
            w190=> c0_n21_w190, 
            w191=> c0_n21_w191, 
            w192=> c0_n21_w192, 
            w193=> c0_n21_w193, 
            w194=> c0_n21_w194, 
            w195=> c0_n21_w195, 
            w196=> c0_n21_w196, 
            w197=> c0_n21_w197, 
            w198=> c0_n21_w198, 
            w199=> c0_n21_w199, 
            w200=> c0_n21_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n21_y
   );           
            
neuron_inst_22: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n22_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n22_w1, 
            w2=> c0_n22_w2, 
            w3=> c0_n22_w3, 
            w4=> c0_n22_w4, 
            w5=> c0_n22_w5, 
            w6=> c0_n22_w6, 
            w7=> c0_n22_w7, 
            w8=> c0_n22_w8, 
            w9=> c0_n22_w9, 
            w10=> c0_n22_w10, 
            w11=> c0_n22_w11, 
            w12=> c0_n22_w12, 
            w13=> c0_n22_w13, 
            w14=> c0_n22_w14, 
            w15=> c0_n22_w15, 
            w16=> c0_n22_w16, 
            w17=> c0_n22_w17, 
            w18=> c0_n22_w18, 
            w19=> c0_n22_w19, 
            w20=> c0_n22_w20, 
            w21=> c0_n22_w21, 
            w22=> c0_n22_w22, 
            w23=> c0_n22_w23, 
            w24=> c0_n22_w24, 
            w25=> c0_n22_w25, 
            w26=> c0_n22_w26, 
            w27=> c0_n22_w27, 
            w28=> c0_n22_w28, 
            w29=> c0_n22_w29, 
            w30=> c0_n22_w30, 
            w31=> c0_n22_w31, 
            w32=> c0_n22_w32, 
            w33=> c0_n22_w33, 
            w34=> c0_n22_w34, 
            w35=> c0_n22_w35, 
            w36=> c0_n22_w36, 
            w37=> c0_n22_w37, 
            w38=> c0_n22_w38, 
            w39=> c0_n22_w39, 
            w40=> c0_n22_w40, 
            w41=> c0_n22_w41, 
            w42=> c0_n22_w42, 
            w43=> c0_n22_w43, 
            w44=> c0_n22_w44, 
            w45=> c0_n22_w45, 
            w46=> c0_n22_w46, 
            w47=> c0_n22_w47, 
            w48=> c0_n22_w48, 
            w49=> c0_n22_w49, 
            w50=> c0_n22_w50, 
            w51=> c0_n22_w51, 
            w52=> c0_n22_w52, 
            w53=> c0_n22_w53, 
            w54=> c0_n22_w54, 
            w55=> c0_n22_w55, 
            w56=> c0_n22_w56, 
            w57=> c0_n22_w57, 
            w58=> c0_n22_w58, 
            w59=> c0_n22_w59, 
            w60=> c0_n22_w60, 
            w61=> c0_n22_w61, 
            w62=> c0_n22_w62, 
            w63=> c0_n22_w63, 
            w64=> c0_n22_w64, 
            w65=> c0_n22_w65, 
            w66=> c0_n22_w66, 
            w67=> c0_n22_w67, 
            w68=> c0_n22_w68, 
            w69=> c0_n22_w69, 
            w70=> c0_n22_w70, 
            w71=> c0_n22_w71, 
            w72=> c0_n22_w72, 
            w73=> c0_n22_w73, 
            w74=> c0_n22_w74, 
            w75=> c0_n22_w75, 
            w76=> c0_n22_w76, 
            w77=> c0_n22_w77, 
            w78=> c0_n22_w78, 
            w79=> c0_n22_w79, 
            w80=> c0_n22_w80, 
            w81=> c0_n22_w81, 
            w82=> c0_n22_w82, 
            w83=> c0_n22_w83, 
            w84=> c0_n22_w84, 
            w85=> c0_n22_w85, 
            w86=> c0_n22_w86, 
            w87=> c0_n22_w87, 
            w88=> c0_n22_w88, 
            w89=> c0_n22_w89, 
            w90=> c0_n22_w90, 
            w91=> c0_n22_w91, 
            w92=> c0_n22_w92, 
            w93=> c0_n22_w93, 
            w94=> c0_n22_w94, 
            w95=> c0_n22_w95, 
            w96=> c0_n22_w96, 
            w97=> c0_n22_w97, 
            w98=> c0_n22_w98, 
            w99=> c0_n22_w99, 
            w100=> c0_n22_w100, 
            w101=> c0_n22_w101, 
            w102=> c0_n22_w102, 
            w103=> c0_n22_w103, 
            w104=> c0_n22_w104, 
            w105=> c0_n22_w105, 
            w106=> c0_n22_w106, 
            w107=> c0_n22_w107, 
            w108=> c0_n22_w108, 
            w109=> c0_n22_w109, 
            w110=> c0_n22_w110, 
            w111=> c0_n22_w111, 
            w112=> c0_n22_w112, 
            w113=> c0_n22_w113, 
            w114=> c0_n22_w114, 
            w115=> c0_n22_w115, 
            w116=> c0_n22_w116, 
            w117=> c0_n22_w117, 
            w118=> c0_n22_w118, 
            w119=> c0_n22_w119, 
            w120=> c0_n22_w120, 
            w121=> c0_n22_w121, 
            w122=> c0_n22_w122, 
            w123=> c0_n22_w123, 
            w124=> c0_n22_w124, 
            w125=> c0_n22_w125, 
            w126=> c0_n22_w126, 
            w127=> c0_n22_w127, 
            w128=> c0_n22_w128, 
            w129=> c0_n22_w129, 
            w130=> c0_n22_w130, 
            w131=> c0_n22_w131, 
            w132=> c0_n22_w132, 
            w133=> c0_n22_w133, 
            w134=> c0_n22_w134, 
            w135=> c0_n22_w135, 
            w136=> c0_n22_w136, 
            w137=> c0_n22_w137, 
            w138=> c0_n22_w138, 
            w139=> c0_n22_w139, 
            w140=> c0_n22_w140, 
            w141=> c0_n22_w141, 
            w142=> c0_n22_w142, 
            w143=> c0_n22_w143, 
            w144=> c0_n22_w144, 
            w145=> c0_n22_w145, 
            w146=> c0_n22_w146, 
            w147=> c0_n22_w147, 
            w148=> c0_n22_w148, 
            w149=> c0_n22_w149, 
            w150=> c0_n22_w150, 
            w151=> c0_n22_w151, 
            w152=> c0_n22_w152, 
            w153=> c0_n22_w153, 
            w154=> c0_n22_w154, 
            w155=> c0_n22_w155, 
            w156=> c0_n22_w156, 
            w157=> c0_n22_w157, 
            w158=> c0_n22_w158, 
            w159=> c0_n22_w159, 
            w160=> c0_n22_w160, 
            w161=> c0_n22_w161, 
            w162=> c0_n22_w162, 
            w163=> c0_n22_w163, 
            w164=> c0_n22_w164, 
            w165=> c0_n22_w165, 
            w166=> c0_n22_w166, 
            w167=> c0_n22_w167, 
            w168=> c0_n22_w168, 
            w169=> c0_n22_w169, 
            w170=> c0_n22_w170, 
            w171=> c0_n22_w171, 
            w172=> c0_n22_w172, 
            w173=> c0_n22_w173, 
            w174=> c0_n22_w174, 
            w175=> c0_n22_w175, 
            w176=> c0_n22_w176, 
            w177=> c0_n22_w177, 
            w178=> c0_n22_w178, 
            w179=> c0_n22_w179, 
            w180=> c0_n22_w180, 
            w181=> c0_n22_w181, 
            w182=> c0_n22_w182, 
            w183=> c0_n22_w183, 
            w184=> c0_n22_w184, 
            w185=> c0_n22_w185, 
            w186=> c0_n22_w186, 
            w187=> c0_n22_w187, 
            w188=> c0_n22_w188, 
            w189=> c0_n22_w189, 
            w190=> c0_n22_w190, 
            w191=> c0_n22_w191, 
            w192=> c0_n22_w192, 
            w193=> c0_n22_w193, 
            w194=> c0_n22_w194, 
            w195=> c0_n22_w195, 
            w196=> c0_n22_w196, 
            w197=> c0_n22_w197, 
            w198=> c0_n22_w198, 
            w199=> c0_n22_w199, 
            w200=> c0_n22_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n22_y
   );           
            
neuron_inst_23: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n23_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n23_w1, 
            w2=> c0_n23_w2, 
            w3=> c0_n23_w3, 
            w4=> c0_n23_w4, 
            w5=> c0_n23_w5, 
            w6=> c0_n23_w6, 
            w7=> c0_n23_w7, 
            w8=> c0_n23_w8, 
            w9=> c0_n23_w9, 
            w10=> c0_n23_w10, 
            w11=> c0_n23_w11, 
            w12=> c0_n23_w12, 
            w13=> c0_n23_w13, 
            w14=> c0_n23_w14, 
            w15=> c0_n23_w15, 
            w16=> c0_n23_w16, 
            w17=> c0_n23_w17, 
            w18=> c0_n23_w18, 
            w19=> c0_n23_w19, 
            w20=> c0_n23_w20, 
            w21=> c0_n23_w21, 
            w22=> c0_n23_w22, 
            w23=> c0_n23_w23, 
            w24=> c0_n23_w24, 
            w25=> c0_n23_w25, 
            w26=> c0_n23_w26, 
            w27=> c0_n23_w27, 
            w28=> c0_n23_w28, 
            w29=> c0_n23_w29, 
            w30=> c0_n23_w30, 
            w31=> c0_n23_w31, 
            w32=> c0_n23_w32, 
            w33=> c0_n23_w33, 
            w34=> c0_n23_w34, 
            w35=> c0_n23_w35, 
            w36=> c0_n23_w36, 
            w37=> c0_n23_w37, 
            w38=> c0_n23_w38, 
            w39=> c0_n23_w39, 
            w40=> c0_n23_w40, 
            w41=> c0_n23_w41, 
            w42=> c0_n23_w42, 
            w43=> c0_n23_w43, 
            w44=> c0_n23_w44, 
            w45=> c0_n23_w45, 
            w46=> c0_n23_w46, 
            w47=> c0_n23_w47, 
            w48=> c0_n23_w48, 
            w49=> c0_n23_w49, 
            w50=> c0_n23_w50, 
            w51=> c0_n23_w51, 
            w52=> c0_n23_w52, 
            w53=> c0_n23_w53, 
            w54=> c0_n23_w54, 
            w55=> c0_n23_w55, 
            w56=> c0_n23_w56, 
            w57=> c0_n23_w57, 
            w58=> c0_n23_w58, 
            w59=> c0_n23_w59, 
            w60=> c0_n23_w60, 
            w61=> c0_n23_w61, 
            w62=> c0_n23_w62, 
            w63=> c0_n23_w63, 
            w64=> c0_n23_w64, 
            w65=> c0_n23_w65, 
            w66=> c0_n23_w66, 
            w67=> c0_n23_w67, 
            w68=> c0_n23_w68, 
            w69=> c0_n23_w69, 
            w70=> c0_n23_w70, 
            w71=> c0_n23_w71, 
            w72=> c0_n23_w72, 
            w73=> c0_n23_w73, 
            w74=> c0_n23_w74, 
            w75=> c0_n23_w75, 
            w76=> c0_n23_w76, 
            w77=> c0_n23_w77, 
            w78=> c0_n23_w78, 
            w79=> c0_n23_w79, 
            w80=> c0_n23_w80, 
            w81=> c0_n23_w81, 
            w82=> c0_n23_w82, 
            w83=> c0_n23_w83, 
            w84=> c0_n23_w84, 
            w85=> c0_n23_w85, 
            w86=> c0_n23_w86, 
            w87=> c0_n23_w87, 
            w88=> c0_n23_w88, 
            w89=> c0_n23_w89, 
            w90=> c0_n23_w90, 
            w91=> c0_n23_w91, 
            w92=> c0_n23_w92, 
            w93=> c0_n23_w93, 
            w94=> c0_n23_w94, 
            w95=> c0_n23_w95, 
            w96=> c0_n23_w96, 
            w97=> c0_n23_w97, 
            w98=> c0_n23_w98, 
            w99=> c0_n23_w99, 
            w100=> c0_n23_w100, 
            w101=> c0_n23_w101, 
            w102=> c0_n23_w102, 
            w103=> c0_n23_w103, 
            w104=> c0_n23_w104, 
            w105=> c0_n23_w105, 
            w106=> c0_n23_w106, 
            w107=> c0_n23_w107, 
            w108=> c0_n23_w108, 
            w109=> c0_n23_w109, 
            w110=> c0_n23_w110, 
            w111=> c0_n23_w111, 
            w112=> c0_n23_w112, 
            w113=> c0_n23_w113, 
            w114=> c0_n23_w114, 
            w115=> c0_n23_w115, 
            w116=> c0_n23_w116, 
            w117=> c0_n23_w117, 
            w118=> c0_n23_w118, 
            w119=> c0_n23_w119, 
            w120=> c0_n23_w120, 
            w121=> c0_n23_w121, 
            w122=> c0_n23_w122, 
            w123=> c0_n23_w123, 
            w124=> c0_n23_w124, 
            w125=> c0_n23_w125, 
            w126=> c0_n23_w126, 
            w127=> c0_n23_w127, 
            w128=> c0_n23_w128, 
            w129=> c0_n23_w129, 
            w130=> c0_n23_w130, 
            w131=> c0_n23_w131, 
            w132=> c0_n23_w132, 
            w133=> c0_n23_w133, 
            w134=> c0_n23_w134, 
            w135=> c0_n23_w135, 
            w136=> c0_n23_w136, 
            w137=> c0_n23_w137, 
            w138=> c0_n23_w138, 
            w139=> c0_n23_w139, 
            w140=> c0_n23_w140, 
            w141=> c0_n23_w141, 
            w142=> c0_n23_w142, 
            w143=> c0_n23_w143, 
            w144=> c0_n23_w144, 
            w145=> c0_n23_w145, 
            w146=> c0_n23_w146, 
            w147=> c0_n23_w147, 
            w148=> c0_n23_w148, 
            w149=> c0_n23_w149, 
            w150=> c0_n23_w150, 
            w151=> c0_n23_w151, 
            w152=> c0_n23_w152, 
            w153=> c0_n23_w153, 
            w154=> c0_n23_w154, 
            w155=> c0_n23_w155, 
            w156=> c0_n23_w156, 
            w157=> c0_n23_w157, 
            w158=> c0_n23_w158, 
            w159=> c0_n23_w159, 
            w160=> c0_n23_w160, 
            w161=> c0_n23_w161, 
            w162=> c0_n23_w162, 
            w163=> c0_n23_w163, 
            w164=> c0_n23_w164, 
            w165=> c0_n23_w165, 
            w166=> c0_n23_w166, 
            w167=> c0_n23_w167, 
            w168=> c0_n23_w168, 
            w169=> c0_n23_w169, 
            w170=> c0_n23_w170, 
            w171=> c0_n23_w171, 
            w172=> c0_n23_w172, 
            w173=> c0_n23_w173, 
            w174=> c0_n23_w174, 
            w175=> c0_n23_w175, 
            w176=> c0_n23_w176, 
            w177=> c0_n23_w177, 
            w178=> c0_n23_w178, 
            w179=> c0_n23_w179, 
            w180=> c0_n23_w180, 
            w181=> c0_n23_w181, 
            w182=> c0_n23_w182, 
            w183=> c0_n23_w183, 
            w184=> c0_n23_w184, 
            w185=> c0_n23_w185, 
            w186=> c0_n23_w186, 
            w187=> c0_n23_w187, 
            w188=> c0_n23_w188, 
            w189=> c0_n23_w189, 
            w190=> c0_n23_w190, 
            w191=> c0_n23_w191, 
            w192=> c0_n23_w192, 
            w193=> c0_n23_w193, 
            w194=> c0_n23_w194, 
            w195=> c0_n23_w195, 
            w196=> c0_n23_w196, 
            w197=> c0_n23_w197, 
            w198=> c0_n23_w198, 
            w199=> c0_n23_w199, 
            w200=> c0_n23_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n23_y
   );           
            
neuron_inst_24: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n24_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n24_w1, 
            w2=> c0_n24_w2, 
            w3=> c0_n24_w3, 
            w4=> c0_n24_w4, 
            w5=> c0_n24_w5, 
            w6=> c0_n24_w6, 
            w7=> c0_n24_w7, 
            w8=> c0_n24_w8, 
            w9=> c0_n24_w9, 
            w10=> c0_n24_w10, 
            w11=> c0_n24_w11, 
            w12=> c0_n24_w12, 
            w13=> c0_n24_w13, 
            w14=> c0_n24_w14, 
            w15=> c0_n24_w15, 
            w16=> c0_n24_w16, 
            w17=> c0_n24_w17, 
            w18=> c0_n24_w18, 
            w19=> c0_n24_w19, 
            w20=> c0_n24_w20, 
            w21=> c0_n24_w21, 
            w22=> c0_n24_w22, 
            w23=> c0_n24_w23, 
            w24=> c0_n24_w24, 
            w25=> c0_n24_w25, 
            w26=> c0_n24_w26, 
            w27=> c0_n24_w27, 
            w28=> c0_n24_w28, 
            w29=> c0_n24_w29, 
            w30=> c0_n24_w30, 
            w31=> c0_n24_w31, 
            w32=> c0_n24_w32, 
            w33=> c0_n24_w33, 
            w34=> c0_n24_w34, 
            w35=> c0_n24_w35, 
            w36=> c0_n24_w36, 
            w37=> c0_n24_w37, 
            w38=> c0_n24_w38, 
            w39=> c0_n24_w39, 
            w40=> c0_n24_w40, 
            w41=> c0_n24_w41, 
            w42=> c0_n24_w42, 
            w43=> c0_n24_w43, 
            w44=> c0_n24_w44, 
            w45=> c0_n24_w45, 
            w46=> c0_n24_w46, 
            w47=> c0_n24_w47, 
            w48=> c0_n24_w48, 
            w49=> c0_n24_w49, 
            w50=> c0_n24_w50, 
            w51=> c0_n24_w51, 
            w52=> c0_n24_w52, 
            w53=> c0_n24_w53, 
            w54=> c0_n24_w54, 
            w55=> c0_n24_w55, 
            w56=> c0_n24_w56, 
            w57=> c0_n24_w57, 
            w58=> c0_n24_w58, 
            w59=> c0_n24_w59, 
            w60=> c0_n24_w60, 
            w61=> c0_n24_w61, 
            w62=> c0_n24_w62, 
            w63=> c0_n24_w63, 
            w64=> c0_n24_w64, 
            w65=> c0_n24_w65, 
            w66=> c0_n24_w66, 
            w67=> c0_n24_w67, 
            w68=> c0_n24_w68, 
            w69=> c0_n24_w69, 
            w70=> c0_n24_w70, 
            w71=> c0_n24_w71, 
            w72=> c0_n24_w72, 
            w73=> c0_n24_w73, 
            w74=> c0_n24_w74, 
            w75=> c0_n24_w75, 
            w76=> c0_n24_w76, 
            w77=> c0_n24_w77, 
            w78=> c0_n24_w78, 
            w79=> c0_n24_w79, 
            w80=> c0_n24_w80, 
            w81=> c0_n24_w81, 
            w82=> c0_n24_w82, 
            w83=> c0_n24_w83, 
            w84=> c0_n24_w84, 
            w85=> c0_n24_w85, 
            w86=> c0_n24_w86, 
            w87=> c0_n24_w87, 
            w88=> c0_n24_w88, 
            w89=> c0_n24_w89, 
            w90=> c0_n24_w90, 
            w91=> c0_n24_w91, 
            w92=> c0_n24_w92, 
            w93=> c0_n24_w93, 
            w94=> c0_n24_w94, 
            w95=> c0_n24_w95, 
            w96=> c0_n24_w96, 
            w97=> c0_n24_w97, 
            w98=> c0_n24_w98, 
            w99=> c0_n24_w99, 
            w100=> c0_n24_w100, 
            w101=> c0_n24_w101, 
            w102=> c0_n24_w102, 
            w103=> c0_n24_w103, 
            w104=> c0_n24_w104, 
            w105=> c0_n24_w105, 
            w106=> c0_n24_w106, 
            w107=> c0_n24_w107, 
            w108=> c0_n24_w108, 
            w109=> c0_n24_w109, 
            w110=> c0_n24_w110, 
            w111=> c0_n24_w111, 
            w112=> c0_n24_w112, 
            w113=> c0_n24_w113, 
            w114=> c0_n24_w114, 
            w115=> c0_n24_w115, 
            w116=> c0_n24_w116, 
            w117=> c0_n24_w117, 
            w118=> c0_n24_w118, 
            w119=> c0_n24_w119, 
            w120=> c0_n24_w120, 
            w121=> c0_n24_w121, 
            w122=> c0_n24_w122, 
            w123=> c0_n24_w123, 
            w124=> c0_n24_w124, 
            w125=> c0_n24_w125, 
            w126=> c0_n24_w126, 
            w127=> c0_n24_w127, 
            w128=> c0_n24_w128, 
            w129=> c0_n24_w129, 
            w130=> c0_n24_w130, 
            w131=> c0_n24_w131, 
            w132=> c0_n24_w132, 
            w133=> c0_n24_w133, 
            w134=> c0_n24_w134, 
            w135=> c0_n24_w135, 
            w136=> c0_n24_w136, 
            w137=> c0_n24_w137, 
            w138=> c0_n24_w138, 
            w139=> c0_n24_w139, 
            w140=> c0_n24_w140, 
            w141=> c0_n24_w141, 
            w142=> c0_n24_w142, 
            w143=> c0_n24_w143, 
            w144=> c0_n24_w144, 
            w145=> c0_n24_w145, 
            w146=> c0_n24_w146, 
            w147=> c0_n24_w147, 
            w148=> c0_n24_w148, 
            w149=> c0_n24_w149, 
            w150=> c0_n24_w150, 
            w151=> c0_n24_w151, 
            w152=> c0_n24_w152, 
            w153=> c0_n24_w153, 
            w154=> c0_n24_w154, 
            w155=> c0_n24_w155, 
            w156=> c0_n24_w156, 
            w157=> c0_n24_w157, 
            w158=> c0_n24_w158, 
            w159=> c0_n24_w159, 
            w160=> c0_n24_w160, 
            w161=> c0_n24_w161, 
            w162=> c0_n24_w162, 
            w163=> c0_n24_w163, 
            w164=> c0_n24_w164, 
            w165=> c0_n24_w165, 
            w166=> c0_n24_w166, 
            w167=> c0_n24_w167, 
            w168=> c0_n24_w168, 
            w169=> c0_n24_w169, 
            w170=> c0_n24_w170, 
            w171=> c0_n24_w171, 
            w172=> c0_n24_w172, 
            w173=> c0_n24_w173, 
            w174=> c0_n24_w174, 
            w175=> c0_n24_w175, 
            w176=> c0_n24_w176, 
            w177=> c0_n24_w177, 
            w178=> c0_n24_w178, 
            w179=> c0_n24_w179, 
            w180=> c0_n24_w180, 
            w181=> c0_n24_w181, 
            w182=> c0_n24_w182, 
            w183=> c0_n24_w183, 
            w184=> c0_n24_w184, 
            w185=> c0_n24_w185, 
            w186=> c0_n24_w186, 
            w187=> c0_n24_w187, 
            w188=> c0_n24_w188, 
            w189=> c0_n24_w189, 
            w190=> c0_n24_w190, 
            w191=> c0_n24_w191, 
            w192=> c0_n24_w192, 
            w193=> c0_n24_w193, 
            w194=> c0_n24_w194, 
            w195=> c0_n24_w195, 
            w196=> c0_n24_w196, 
            w197=> c0_n24_w197, 
            w198=> c0_n24_w198, 
            w199=> c0_n24_w199, 
            w200=> c0_n24_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n24_y
   );           
            
neuron_inst_25: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n25_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n25_w1, 
            w2=> c0_n25_w2, 
            w3=> c0_n25_w3, 
            w4=> c0_n25_w4, 
            w5=> c0_n25_w5, 
            w6=> c0_n25_w6, 
            w7=> c0_n25_w7, 
            w8=> c0_n25_w8, 
            w9=> c0_n25_w9, 
            w10=> c0_n25_w10, 
            w11=> c0_n25_w11, 
            w12=> c0_n25_w12, 
            w13=> c0_n25_w13, 
            w14=> c0_n25_w14, 
            w15=> c0_n25_w15, 
            w16=> c0_n25_w16, 
            w17=> c0_n25_w17, 
            w18=> c0_n25_w18, 
            w19=> c0_n25_w19, 
            w20=> c0_n25_w20, 
            w21=> c0_n25_w21, 
            w22=> c0_n25_w22, 
            w23=> c0_n25_w23, 
            w24=> c0_n25_w24, 
            w25=> c0_n25_w25, 
            w26=> c0_n25_w26, 
            w27=> c0_n25_w27, 
            w28=> c0_n25_w28, 
            w29=> c0_n25_w29, 
            w30=> c0_n25_w30, 
            w31=> c0_n25_w31, 
            w32=> c0_n25_w32, 
            w33=> c0_n25_w33, 
            w34=> c0_n25_w34, 
            w35=> c0_n25_w35, 
            w36=> c0_n25_w36, 
            w37=> c0_n25_w37, 
            w38=> c0_n25_w38, 
            w39=> c0_n25_w39, 
            w40=> c0_n25_w40, 
            w41=> c0_n25_w41, 
            w42=> c0_n25_w42, 
            w43=> c0_n25_w43, 
            w44=> c0_n25_w44, 
            w45=> c0_n25_w45, 
            w46=> c0_n25_w46, 
            w47=> c0_n25_w47, 
            w48=> c0_n25_w48, 
            w49=> c0_n25_w49, 
            w50=> c0_n25_w50, 
            w51=> c0_n25_w51, 
            w52=> c0_n25_w52, 
            w53=> c0_n25_w53, 
            w54=> c0_n25_w54, 
            w55=> c0_n25_w55, 
            w56=> c0_n25_w56, 
            w57=> c0_n25_w57, 
            w58=> c0_n25_w58, 
            w59=> c0_n25_w59, 
            w60=> c0_n25_w60, 
            w61=> c0_n25_w61, 
            w62=> c0_n25_w62, 
            w63=> c0_n25_w63, 
            w64=> c0_n25_w64, 
            w65=> c0_n25_w65, 
            w66=> c0_n25_w66, 
            w67=> c0_n25_w67, 
            w68=> c0_n25_w68, 
            w69=> c0_n25_w69, 
            w70=> c0_n25_w70, 
            w71=> c0_n25_w71, 
            w72=> c0_n25_w72, 
            w73=> c0_n25_w73, 
            w74=> c0_n25_w74, 
            w75=> c0_n25_w75, 
            w76=> c0_n25_w76, 
            w77=> c0_n25_w77, 
            w78=> c0_n25_w78, 
            w79=> c0_n25_w79, 
            w80=> c0_n25_w80, 
            w81=> c0_n25_w81, 
            w82=> c0_n25_w82, 
            w83=> c0_n25_w83, 
            w84=> c0_n25_w84, 
            w85=> c0_n25_w85, 
            w86=> c0_n25_w86, 
            w87=> c0_n25_w87, 
            w88=> c0_n25_w88, 
            w89=> c0_n25_w89, 
            w90=> c0_n25_w90, 
            w91=> c0_n25_w91, 
            w92=> c0_n25_w92, 
            w93=> c0_n25_w93, 
            w94=> c0_n25_w94, 
            w95=> c0_n25_w95, 
            w96=> c0_n25_w96, 
            w97=> c0_n25_w97, 
            w98=> c0_n25_w98, 
            w99=> c0_n25_w99, 
            w100=> c0_n25_w100, 
            w101=> c0_n25_w101, 
            w102=> c0_n25_w102, 
            w103=> c0_n25_w103, 
            w104=> c0_n25_w104, 
            w105=> c0_n25_w105, 
            w106=> c0_n25_w106, 
            w107=> c0_n25_w107, 
            w108=> c0_n25_w108, 
            w109=> c0_n25_w109, 
            w110=> c0_n25_w110, 
            w111=> c0_n25_w111, 
            w112=> c0_n25_w112, 
            w113=> c0_n25_w113, 
            w114=> c0_n25_w114, 
            w115=> c0_n25_w115, 
            w116=> c0_n25_w116, 
            w117=> c0_n25_w117, 
            w118=> c0_n25_w118, 
            w119=> c0_n25_w119, 
            w120=> c0_n25_w120, 
            w121=> c0_n25_w121, 
            w122=> c0_n25_w122, 
            w123=> c0_n25_w123, 
            w124=> c0_n25_w124, 
            w125=> c0_n25_w125, 
            w126=> c0_n25_w126, 
            w127=> c0_n25_w127, 
            w128=> c0_n25_w128, 
            w129=> c0_n25_w129, 
            w130=> c0_n25_w130, 
            w131=> c0_n25_w131, 
            w132=> c0_n25_w132, 
            w133=> c0_n25_w133, 
            w134=> c0_n25_w134, 
            w135=> c0_n25_w135, 
            w136=> c0_n25_w136, 
            w137=> c0_n25_w137, 
            w138=> c0_n25_w138, 
            w139=> c0_n25_w139, 
            w140=> c0_n25_w140, 
            w141=> c0_n25_w141, 
            w142=> c0_n25_w142, 
            w143=> c0_n25_w143, 
            w144=> c0_n25_w144, 
            w145=> c0_n25_w145, 
            w146=> c0_n25_w146, 
            w147=> c0_n25_w147, 
            w148=> c0_n25_w148, 
            w149=> c0_n25_w149, 
            w150=> c0_n25_w150, 
            w151=> c0_n25_w151, 
            w152=> c0_n25_w152, 
            w153=> c0_n25_w153, 
            w154=> c0_n25_w154, 
            w155=> c0_n25_w155, 
            w156=> c0_n25_w156, 
            w157=> c0_n25_w157, 
            w158=> c0_n25_w158, 
            w159=> c0_n25_w159, 
            w160=> c0_n25_w160, 
            w161=> c0_n25_w161, 
            w162=> c0_n25_w162, 
            w163=> c0_n25_w163, 
            w164=> c0_n25_w164, 
            w165=> c0_n25_w165, 
            w166=> c0_n25_w166, 
            w167=> c0_n25_w167, 
            w168=> c0_n25_w168, 
            w169=> c0_n25_w169, 
            w170=> c0_n25_w170, 
            w171=> c0_n25_w171, 
            w172=> c0_n25_w172, 
            w173=> c0_n25_w173, 
            w174=> c0_n25_w174, 
            w175=> c0_n25_w175, 
            w176=> c0_n25_w176, 
            w177=> c0_n25_w177, 
            w178=> c0_n25_w178, 
            w179=> c0_n25_w179, 
            w180=> c0_n25_w180, 
            w181=> c0_n25_w181, 
            w182=> c0_n25_w182, 
            w183=> c0_n25_w183, 
            w184=> c0_n25_w184, 
            w185=> c0_n25_w185, 
            w186=> c0_n25_w186, 
            w187=> c0_n25_w187, 
            w188=> c0_n25_w188, 
            w189=> c0_n25_w189, 
            w190=> c0_n25_w190, 
            w191=> c0_n25_w191, 
            w192=> c0_n25_w192, 
            w193=> c0_n25_w193, 
            w194=> c0_n25_w194, 
            w195=> c0_n25_w195, 
            w196=> c0_n25_w196, 
            w197=> c0_n25_w197, 
            w198=> c0_n25_w198, 
            w199=> c0_n25_w199, 
            w200=> c0_n25_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n25_y
   );           
            
neuron_inst_26: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n26_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n26_w1, 
            w2=> c0_n26_w2, 
            w3=> c0_n26_w3, 
            w4=> c0_n26_w4, 
            w5=> c0_n26_w5, 
            w6=> c0_n26_w6, 
            w7=> c0_n26_w7, 
            w8=> c0_n26_w8, 
            w9=> c0_n26_w9, 
            w10=> c0_n26_w10, 
            w11=> c0_n26_w11, 
            w12=> c0_n26_w12, 
            w13=> c0_n26_w13, 
            w14=> c0_n26_w14, 
            w15=> c0_n26_w15, 
            w16=> c0_n26_w16, 
            w17=> c0_n26_w17, 
            w18=> c0_n26_w18, 
            w19=> c0_n26_w19, 
            w20=> c0_n26_w20, 
            w21=> c0_n26_w21, 
            w22=> c0_n26_w22, 
            w23=> c0_n26_w23, 
            w24=> c0_n26_w24, 
            w25=> c0_n26_w25, 
            w26=> c0_n26_w26, 
            w27=> c0_n26_w27, 
            w28=> c0_n26_w28, 
            w29=> c0_n26_w29, 
            w30=> c0_n26_w30, 
            w31=> c0_n26_w31, 
            w32=> c0_n26_w32, 
            w33=> c0_n26_w33, 
            w34=> c0_n26_w34, 
            w35=> c0_n26_w35, 
            w36=> c0_n26_w36, 
            w37=> c0_n26_w37, 
            w38=> c0_n26_w38, 
            w39=> c0_n26_w39, 
            w40=> c0_n26_w40, 
            w41=> c0_n26_w41, 
            w42=> c0_n26_w42, 
            w43=> c0_n26_w43, 
            w44=> c0_n26_w44, 
            w45=> c0_n26_w45, 
            w46=> c0_n26_w46, 
            w47=> c0_n26_w47, 
            w48=> c0_n26_w48, 
            w49=> c0_n26_w49, 
            w50=> c0_n26_w50, 
            w51=> c0_n26_w51, 
            w52=> c0_n26_w52, 
            w53=> c0_n26_w53, 
            w54=> c0_n26_w54, 
            w55=> c0_n26_w55, 
            w56=> c0_n26_w56, 
            w57=> c0_n26_w57, 
            w58=> c0_n26_w58, 
            w59=> c0_n26_w59, 
            w60=> c0_n26_w60, 
            w61=> c0_n26_w61, 
            w62=> c0_n26_w62, 
            w63=> c0_n26_w63, 
            w64=> c0_n26_w64, 
            w65=> c0_n26_w65, 
            w66=> c0_n26_w66, 
            w67=> c0_n26_w67, 
            w68=> c0_n26_w68, 
            w69=> c0_n26_w69, 
            w70=> c0_n26_w70, 
            w71=> c0_n26_w71, 
            w72=> c0_n26_w72, 
            w73=> c0_n26_w73, 
            w74=> c0_n26_w74, 
            w75=> c0_n26_w75, 
            w76=> c0_n26_w76, 
            w77=> c0_n26_w77, 
            w78=> c0_n26_w78, 
            w79=> c0_n26_w79, 
            w80=> c0_n26_w80, 
            w81=> c0_n26_w81, 
            w82=> c0_n26_w82, 
            w83=> c0_n26_w83, 
            w84=> c0_n26_w84, 
            w85=> c0_n26_w85, 
            w86=> c0_n26_w86, 
            w87=> c0_n26_w87, 
            w88=> c0_n26_w88, 
            w89=> c0_n26_w89, 
            w90=> c0_n26_w90, 
            w91=> c0_n26_w91, 
            w92=> c0_n26_w92, 
            w93=> c0_n26_w93, 
            w94=> c0_n26_w94, 
            w95=> c0_n26_w95, 
            w96=> c0_n26_w96, 
            w97=> c0_n26_w97, 
            w98=> c0_n26_w98, 
            w99=> c0_n26_w99, 
            w100=> c0_n26_w100, 
            w101=> c0_n26_w101, 
            w102=> c0_n26_w102, 
            w103=> c0_n26_w103, 
            w104=> c0_n26_w104, 
            w105=> c0_n26_w105, 
            w106=> c0_n26_w106, 
            w107=> c0_n26_w107, 
            w108=> c0_n26_w108, 
            w109=> c0_n26_w109, 
            w110=> c0_n26_w110, 
            w111=> c0_n26_w111, 
            w112=> c0_n26_w112, 
            w113=> c0_n26_w113, 
            w114=> c0_n26_w114, 
            w115=> c0_n26_w115, 
            w116=> c0_n26_w116, 
            w117=> c0_n26_w117, 
            w118=> c0_n26_w118, 
            w119=> c0_n26_w119, 
            w120=> c0_n26_w120, 
            w121=> c0_n26_w121, 
            w122=> c0_n26_w122, 
            w123=> c0_n26_w123, 
            w124=> c0_n26_w124, 
            w125=> c0_n26_w125, 
            w126=> c0_n26_w126, 
            w127=> c0_n26_w127, 
            w128=> c0_n26_w128, 
            w129=> c0_n26_w129, 
            w130=> c0_n26_w130, 
            w131=> c0_n26_w131, 
            w132=> c0_n26_w132, 
            w133=> c0_n26_w133, 
            w134=> c0_n26_w134, 
            w135=> c0_n26_w135, 
            w136=> c0_n26_w136, 
            w137=> c0_n26_w137, 
            w138=> c0_n26_w138, 
            w139=> c0_n26_w139, 
            w140=> c0_n26_w140, 
            w141=> c0_n26_w141, 
            w142=> c0_n26_w142, 
            w143=> c0_n26_w143, 
            w144=> c0_n26_w144, 
            w145=> c0_n26_w145, 
            w146=> c0_n26_w146, 
            w147=> c0_n26_w147, 
            w148=> c0_n26_w148, 
            w149=> c0_n26_w149, 
            w150=> c0_n26_w150, 
            w151=> c0_n26_w151, 
            w152=> c0_n26_w152, 
            w153=> c0_n26_w153, 
            w154=> c0_n26_w154, 
            w155=> c0_n26_w155, 
            w156=> c0_n26_w156, 
            w157=> c0_n26_w157, 
            w158=> c0_n26_w158, 
            w159=> c0_n26_w159, 
            w160=> c0_n26_w160, 
            w161=> c0_n26_w161, 
            w162=> c0_n26_w162, 
            w163=> c0_n26_w163, 
            w164=> c0_n26_w164, 
            w165=> c0_n26_w165, 
            w166=> c0_n26_w166, 
            w167=> c0_n26_w167, 
            w168=> c0_n26_w168, 
            w169=> c0_n26_w169, 
            w170=> c0_n26_w170, 
            w171=> c0_n26_w171, 
            w172=> c0_n26_w172, 
            w173=> c0_n26_w173, 
            w174=> c0_n26_w174, 
            w175=> c0_n26_w175, 
            w176=> c0_n26_w176, 
            w177=> c0_n26_w177, 
            w178=> c0_n26_w178, 
            w179=> c0_n26_w179, 
            w180=> c0_n26_w180, 
            w181=> c0_n26_w181, 
            w182=> c0_n26_w182, 
            w183=> c0_n26_w183, 
            w184=> c0_n26_w184, 
            w185=> c0_n26_w185, 
            w186=> c0_n26_w186, 
            w187=> c0_n26_w187, 
            w188=> c0_n26_w188, 
            w189=> c0_n26_w189, 
            w190=> c0_n26_w190, 
            w191=> c0_n26_w191, 
            w192=> c0_n26_w192, 
            w193=> c0_n26_w193, 
            w194=> c0_n26_w194, 
            w195=> c0_n26_w195, 
            w196=> c0_n26_w196, 
            w197=> c0_n26_w197, 
            w198=> c0_n26_w198, 
            w199=> c0_n26_w199, 
            w200=> c0_n26_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n26_y
   );           
            
neuron_inst_27: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n27_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n27_w1, 
            w2=> c0_n27_w2, 
            w3=> c0_n27_w3, 
            w4=> c0_n27_w4, 
            w5=> c0_n27_w5, 
            w6=> c0_n27_w6, 
            w7=> c0_n27_w7, 
            w8=> c0_n27_w8, 
            w9=> c0_n27_w9, 
            w10=> c0_n27_w10, 
            w11=> c0_n27_w11, 
            w12=> c0_n27_w12, 
            w13=> c0_n27_w13, 
            w14=> c0_n27_w14, 
            w15=> c0_n27_w15, 
            w16=> c0_n27_w16, 
            w17=> c0_n27_w17, 
            w18=> c0_n27_w18, 
            w19=> c0_n27_w19, 
            w20=> c0_n27_w20, 
            w21=> c0_n27_w21, 
            w22=> c0_n27_w22, 
            w23=> c0_n27_w23, 
            w24=> c0_n27_w24, 
            w25=> c0_n27_w25, 
            w26=> c0_n27_w26, 
            w27=> c0_n27_w27, 
            w28=> c0_n27_w28, 
            w29=> c0_n27_w29, 
            w30=> c0_n27_w30, 
            w31=> c0_n27_w31, 
            w32=> c0_n27_w32, 
            w33=> c0_n27_w33, 
            w34=> c0_n27_w34, 
            w35=> c0_n27_w35, 
            w36=> c0_n27_w36, 
            w37=> c0_n27_w37, 
            w38=> c0_n27_w38, 
            w39=> c0_n27_w39, 
            w40=> c0_n27_w40, 
            w41=> c0_n27_w41, 
            w42=> c0_n27_w42, 
            w43=> c0_n27_w43, 
            w44=> c0_n27_w44, 
            w45=> c0_n27_w45, 
            w46=> c0_n27_w46, 
            w47=> c0_n27_w47, 
            w48=> c0_n27_w48, 
            w49=> c0_n27_w49, 
            w50=> c0_n27_w50, 
            w51=> c0_n27_w51, 
            w52=> c0_n27_w52, 
            w53=> c0_n27_w53, 
            w54=> c0_n27_w54, 
            w55=> c0_n27_w55, 
            w56=> c0_n27_w56, 
            w57=> c0_n27_w57, 
            w58=> c0_n27_w58, 
            w59=> c0_n27_w59, 
            w60=> c0_n27_w60, 
            w61=> c0_n27_w61, 
            w62=> c0_n27_w62, 
            w63=> c0_n27_w63, 
            w64=> c0_n27_w64, 
            w65=> c0_n27_w65, 
            w66=> c0_n27_w66, 
            w67=> c0_n27_w67, 
            w68=> c0_n27_w68, 
            w69=> c0_n27_w69, 
            w70=> c0_n27_w70, 
            w71=> c0_n27_w71, 
            w72=> c0_n27_w72, 
            w73=> c0_n27_w73, 
            w74=> c0_n27_w74, 
            w75=> c0_n27_w75, 
            w76=> c0_n27_w76, 
            w77=> c0_n27_w77, 
            w78=> c0_n27_w78, 
            w79=> c0_n27_w79, 
            w80=> c0_n27_w80, 
            w81=> c0_n27_w81, 
            w82=> c0_n27_w82, 
            w83=> c0_n27_w83, 
            w84=> c0_n27_w84, 
            w85=> c0_n27_w85, 
            w86=> c0_n27_w86, 
            w87=> c0_n27_w87, 
            w88=> c0_n27_w88, 
            w89=> c0_n27_w89, 
            w90=> c0_n27_w90, 
            w91=> c0_n27_w91, 
            w92=> c0_n27_w92, 
            w93=> c0_n27_w93, 
            w94=> c0_n27_w94, 
            w95=> c0_n27_w95, 
            w96=> c0_n27_w96, 
            w97=> c0_n27_w97, 
            w98=> c0_n27_w98, 
            w99=> c0_n27_w99, 
            w100=> c0_n27_w100, 
            w101=> c0_n27_w101, 
            w102=> c0_n27_w102, 
            w103=> c0_n27_w103, 
            w104=> c0_n27_w104, 
            w105=> c0_n27_w105, 
            w106=> c0_n27_w106, 
            w107=> c0_n27_w107, 
            w108=> c0_n27_w108, 
            w109=> c0_n27_w109, 
            w110=> c0_n27_w110, 
            w111=> c0_n27_w111, 
            w112=> c0_n27_w112, 
            w113=> c0_n27_w113, 
            w114=> c0_n27_w114, 
            w115=> c0_n27_w115, 
            w116=> c0_n27_w116, 
            w117=> c0_n27_w117, 
            w118=> c0_n27_w118, 
            w119=> c0_n27_w119, 
            w120=> c0_n27_w120, 
            w121=> c0_n27_w121, 
            w122=> c0_n27_w122, 
            w123=> c0_n27_w123, 
            w124=> c0_n27_w124, 
            w125=> c0_n27_w125, 
            w126=> c0_n27_w126, 
            w127=> c0_n27_w127, 
            w128=> c0_n27_w128, 
            w129=> c0_n27_w129, 
            w130=> c0_n27_w130, 
            w131=> c0_n27_w131, 
            w132=> c0_n27_w132, 
            w133=> c0_n27_w133, 
            w134=> c0_n27_w134, 
            w135=> c0_n27_w135, 
            w136=> c0_n27_w136, 
            w137=> c0_n27_w137, 
            w138=> c0_n27_w138, 
            w139=> c0_n27_w139, 
            w140=> c0_n27_w140, 
            w141=> c0_n27_w141, 
            w142=> c0_n27_w142, 
            w143=> c0_n27_w143, 
            w144=> c0_n27_w144, 
            w145=> c0_n27_w145, 
            w146=> c0_n27_w146, 
            w147=> c0_n27_w147, 
            w148=> c0_n27_w148, 
            w149=> c0_n27_w149, 
            w150=> c0_n27_w150, 
            w151=> c0_n27_w151, 
            w152=> c0_n27_w152, 
            w153=> c0_n27_w153, 
            w154=> c0_n27_w154, 
            w155=> c0_n27_w155, 
            w156=> c0_n27_w156, 
            w157=> c0_n27_w157, 
            w158=> c0_n27_w158, 
            w159=> c0_n27_w159, 
            w160=> c0_n27_w160, 
            w161=> c0_n27_w161, 
            w162=> c0_n27_w162, 
            w163=> c0_n27_w163, 
            w164=> c0_n27_w164, 
            w165=> c0_n27_w165, 
            w166=> c0_n27_w166, 
            w167=> c0_n27_w167, 
            w168=> c0_n27_w168, 
            w169=> c0_n27_w169, 
            w170=> c0_n27_w170, 
            w171=> c0_n27_w171, 
            w172=> c0_n27_w172, 
            w173=> c0_n27_w173, 
            w174=> c0_n27_w174, 
            w175=> c0_n27_w175, 
            w176=> c0_n27_w176, 
            w177=> c0_n27_w177, 
            w178=> c0_n27_w178, 
            w179=> c0_n27_w179, 
            w180=> c0_n27_w180, 
            w181=> c0_n27_w181, 
            w182=> c0_n27_w182, 
            w183=> c0_n27_w183, 
            w184=> c0_n27_w184, 
            w185=> c0_n27_w185, 
            w186=> c0_n27_w186, 
            w187=> c0_n27_w187, 
            w188=> c0_n27_w188, 
            w189=> c0_n27_w189, 
            w190=> c0_n27_w190, 
            w191=> c0_n27_w191, 
            w192=> c0_n27_w192, 
            w193=> c0_n27_w193, 
            w194=> c0_n27_w194, 
            w195=> c0_n27_w195, 
            w196=> c0_n27_w196, 
            w197=> c0_n27_w197, 
            w198=> c0_n27_w198, 
            w199=> c0_n27_w199, 
            w200=> c0_n27_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n27_y
   );           
            
neuron_inst_28: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n28_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n28_w1, 
            w2=> c0_n28_w2, 
            w3=> c0_n28_w3, 
            w4=> c0_n28_w4, 
            w5=> c0_n28_w5, 
            w6=> c0_n28_w6, 
            w7=> c0_n28_w7, 
            w8=> c0_n28_w8, 
            w9=> c0_n28_w9, 
            w10=> c0_n28_w10, 
            w11=> c0_n28_w11, 
            w12=> c0_n28_w12, 
            w13=> c0_n28_w13, 
            w14=> c0_n28_w14, 
            w15=> c0_n28_w15, 
            w16=> c0_n28_w16, 
            w17=> c0_n28_w17, 
            w18=> c0_n28_w18, 
            w19=> c0_n28_w19, 
            w20=> c0_n28_w20, 
            w21=> c0_n28_w21, 
            w22=> c0_n28_w22, 
            w23=> c0_n28_w23, 
            w24=> c0_n28_w24, 
            w25=> c0_n28_w25, 
            w26=> c0_n28_w26, 
            w27=> c0_n28_w27, 
            w28=> c0_n28_w28, 
            w29=> c0_n28_w29, 
            w30=> c0_n28_w30, 
            w31=> c0_n28_w31, 
            w32=> c0_n28_w32, 
            w33=> c0_n28_w33, 
            w34=> c0_n28_w34, 
            w35=> c0_n28_w35, 
            w36=> c0_n28_w36, 
            w37=> c0_n28_w37, 
            w38=> c0_n28_w38, 
            w39=> c0_n28_w39, 
            w40=> c0_n28_w40, 
            w41=> c0_n28_w41, 
            w42=> c0_n28_w42, 
            w43=> c0_n28_w43, 
            w44=> c0_n28_w44, 
            w45=> c0_n28_w45, 
            w46=> c0_n28_w46, 
            w47=> c0_n28_w47, 
            w48=> c0_n28_w48, 
            w49=> c0_n28_w49, 
            w50=> c0_n28_w50, 
            w51=> c0_n28_w51, 
            w52=> c0_n28_w52, 
            w53=> c0_n28_w53, 
            w54=> c0_n28_w54, 
            w55=> c0_n28_w55, 
            w56=> c0_n28_w56, 
            w57=> c0_n28_w57, 
            w58=> c0_n28_w58, 
            w59=> c0_n28_w59, 
            w60=> c0_n28_w60, 
            w61=> c0_n28_w61, 
            w62=> c0_n28_w62, 
            w63=> c0_n28_w63, 
            w64=> c0_n28_w64, 
            w65=> c0_n28_w65, 
            w66=> c0_n28_w66, 
            w67=> c0_n28_w67, 
            w68=> c0_n28_w68, 
            w69=> c0_n28_w69, 
            w70=> c0_n28_w70, 
            w71=> c0_n28_w71, 
            w72=> c0_n28_w72, 
            w73=> c0_n28_w73, 
            w74=> c0_n28_w74, 
            w75=> c0_n28_w75, 
            w76=> c0_n28_w76, 
            w77=> c0_n28_w77, 
            w78=> c0_n28_w78, 
            w79=> c0_n28_w79, 
            w80=> c0_n28_w80, 
            w81=> c0_n28_w81, 
            w82=> c0_n28_w82, 
            w83=> c0_n28_w83, 
            w84=> c0_n28_w84, 
            w85=> c0_n28_w85, 
            w86=> c0_n28_w86, 
            w87=> c0_n28_w87, 
            w88=> c0_n28_w88, 
            w89=> c0_n28_w89, 
            w90=> c0_n28_w90, 
            w91=> c0_n28_w91, 
            w92=> c0_n28_w92, 
            w93=> c0_n28_w93, 
            w94=> c0_n28_w94, 
            w95=> c0_n28_w95, 
            w96=> c0_n28_w96, 
            w97=> c0_n28_w97, 
            w98=> c0_n28_w98, 
            w99=> c0_n28_w99, 
            w100=> c0_n28_w100, 
            w101=> c0_n28_w101, 
            w102=> c0_n28_w102, 
            w103=> c0_n28_w103, 
            w104=> c0_n28_w104, 
            w105=> c0_n28_w105, 
            w106=> c0_n28_w106, 
            w107=> c0_n28_w107, 
            w108=> c0_n28_w108, 
            w109=> c0_n28_w109, 
            w110=> c0_n28_w110, 
            w111=> c0_n28_w111, 
            w112=> c0_n28_w112, 
            w113=> c0_n28_w113, 
            w114=> c0_n28_w114, 
            w115=> c0_n28_w115, 
            w116=> c0_n28_w116, 
            w117=> c0_n28_w117, 
            w118=> c0_n28_w118, 
            w119=> c0_n28_w119, 
            w120=> c0_n28_w120, 
            w121=> c0_n28_w121, 
            w122=> c0_n28_w122, 
            w123=> c0_n28_w123, 
            w124=> c0_n28_w124, 
            w125=> c0_n28_w125, 
            w126=> c0_n28_w126, 
            w127=> c0_n28_w127, 
            w128=> c0_n28_w128, 
            w129=> c0_n28_w129, 
            w130=> c0_n28_w130, 
            w131=> c0_n28_w131, 
            w132=> c0_n28_w132, 
            w133=> c0_n28_w133, 
            w134=> c0_n28_w134, 
            w135=> c0_n28_w135, 
            w136=> c0_n28_w136, 
            w137=> c0_n28_w137, 
            w138=> c0_n28_w138, 
            w139=> c0_n28_w139, 
            w140=> c0_n28_w140, 
            w141=> c0_n28_w141, 
            w142=> c0_n28_w142, 
            w143=> c0_n28_w143, 
            w144=> c0_n28_w144, 
            w145=> c0_n28_w145, 
            w146=> c0_n28_w146, 
            w147=> c0_n28_w147, 
            w148=> c0_n28_w148, 
            w149=> c0_n28_w149, 
            w150=> c0_n28_w150, 
            w151=> c0_n28_w151, 
            w152=> c0_n28_w152, 
            w153=> c0_n28_w153, 
            w154=> c0_n28_w154, 
            w155=> c0_n28_w155, 
            w156=> c0_n28_w156, 
            w157=> c0_n28_w157, 
            w158=> c0_n28_w158, 
            w159=> c0_n28_w159, 
            w160=> c0_n28_w160, 
            w161=> c0_n28_w161, 
            w162=> c0_n28_w162, 
            w163=> c0_n28_w163, 
            w164=> c0_n28_w164, 
            w165=> c0_n28_w165, 
            w166=> c0_n28_w166, 
            w167=> c0_n28_w167, 
            w168=> c0_n28_w168, 
            w169=> c0_n28_w169, 
            w170=> c0_n28_w170, 
            w171=> c0_n28_w171, 
            w172=> c0_n28_w172, 
            w173=> c0_n28_w173, 
            w174=> c0_n28_w174, 
            w175=> c0_n28_w175, 
            w176=> c0_n28_w176, 
            w177=> c0_n28_w177, 
            w178=> c0_n28_w178, 
            w179=> c0_n28_w179, 
            w180=> c0_n28_w180, 
            w181=> c0_n28_w181, 
            w182=> c0_n28_w182, 
            w183=> c0_n28_w183, 
            w184=> c0_n28_w184, 
            w185=> c0_n28_w185, 
            w186=> c0_n28_w186, 
            w187=> c0_n28_w187, 
            w188=> c0_n28_w188, 
            w189=> c0_n28_w189, 
            w190=> c0_n28_w190, 
            w191=> c0_n28_w191, 
            w192=> c0_n28_w192, 
            w193=> c0_n28_w193, 
            w194=> c0_n28_w194, 
            w195=> c0_n28_w195, 
            w196=> c0_n28_w196, 
            w197=> c0_n28_w197, 
            w198=> c0_n28_w198, 
            w199=> c0_n28_w199, 
            w200=> c0_n28_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n28_y
   );           
            
neuron_inst_29: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n29_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n29_w1, 
            w2=> c0_n29_w2, 
            w3=> c0_n29_w3, 
            w4=> c0_n29_w4, 
            w5=> c0_n29_w5, 
            w6=> c0_n29_w6, 
            w7=> c0_n29_w7, 
            w8=> c0_n29_w8, 
            w9=> c0_n29_w9, 
            w10=> c0_n29_w10, 
            w11=> c0_n29_w11, 
            w12=> c0_n29_w12, 
            w13=> c0_n29_w13, 
            w14=> c0_n29_w14, 
            w15=> c0_n29_w15, 
            w16=> c0_n29_w16, 
            w17=> c0_n29_w17, 
            w18=> c0_n29_w18, 
            w19=> c0_n29_w19, 
            w20=> c0_n29_w20, 
            w21=> c0_n29_w21, 
            w22=> c0_n29_w22, 
            w23=> c0_n29_w23, 
            w24=> c0_n29_w24, 
            w25=> c0_n29_w25, 
            w26=> c0_n29_w26, 
            w27=> c0_n29_w27, 
            w28=> c0_n29_w28, 
            w29=> c0_n29_w29, 
            w30=> c0_n29_w30, 
            w31=> c0_n29_w31, 
            w32=> c0_n29_w32, 
            w33=> c0_n29_w33, 
            w34=> c0_n29_w34, 
            w35=> c0_n29_w35, 
            w36=> c0_n29_w36, 
            w37=> c0_n29_w37, 
            w38=> c0_n29_w38, 
            w39=> c0_n29_w39, 
            w40=> c0_n29_w40, 
            w41=> c0_n29_w41, 
            w42=> c0_n29_w42, 
            w43=> c0_n29_w43, 
            w44=> c0_n29_w44, 
            w45=> c0_n29_w45, 
            w46=> c0_n29_w46, 
            w47=> c0_n29_w47, 
            w48=> c0_n29_w48, 
            w49=> c0_n29_w49, 
            w50=> c0_n29_w50, 
            w51=> c0_n29_w51, 
            w52=> c0_n29_w52, 
            w53=> c0_n29_w53, 
            w54=> c0_n29_w54, 
            w55=> c0_n29_w55, 
            w56=> c0_n29_w56, 
            w57=> c0_n29_w57, 
            w58=> c0_n29_w58, 
            w59=> c0_n29_w59, 
            w60=> c0_n29_w60, 
            w61=> c0_n29_w61, 
            w62=> c0_n29_w62, 
            w63=> c0_n29_w63, 
            w64=> c0_n29_w64, 
            w65=> c0_n29_w65, 
            w66=> c0_n29_w66, 
            w67=> c0_n29_w67, 
            w68=> c0_n29_w68, 
            w69=> c0_n29_w69, 
            w70=> c0_n29_w70, 
            w71=> c0_n29_w71, 
            w72=> c0_n29_w72, 
            w73=> c0_n29_w73, 
            w74=> c0_n29_w74, 
            w75=> c0_n29_w75, 
            w76=> c0_n29_w76, 
            w77=> c0_n29_w77, 
            w78=> c0_n29_w78, 
            w79=> c0_n29_w79, 
            w80=> c0_n29_w80, 
            w81=> c0_n29_w81, 
            w82=> c0_n29_w82, 
            w83=> c0_n29_w83, 
            w84=> c0_n29_w84, 
            w85=> c0_n29_w85, 
            w86=> c0_n29_w86, 
            w87=> c0_n29_w87, 
            w88=> c0_n29_w88, 
            w89=> c0_n29_w89, 
            w90=> c0_n29_w90, 
            w91=> c0_n29_w91, 
            w92=> c0_n29_w92, 
            w93=> c0_n29_w93, 
            w94=> c0_n29_w94, 
            w95=> c0_n29_w95, 
            w96=> c0_n29_w96, 
            w97=> c0_n29_w97, 
            w98=> c0_n29_w98, 
            w99=> c0_n29_w99, 
            w100=> c0_n29_w100, 
            w101=> c0_n29_w101, 
            w102=> c0_n29_w102, 
            w103=> c0_n29_w103, 
            w104=> c0_n29_w104, 
            w105=> c0_n29_w105, 
            w106=> c0_n29_w106, 
            w107=> c0_n29_w107, 
            w108=> c0_n29_w108, 
            w109=> c0_n29_w109, 
            w110=> c0_n29_w110, 
            w111=> c0_n29_w111, 
            w112=> c0_n29_w112, 
            w113=> c0_n29_w113, 
            w114=> c0_n29_w114, 
            w115=> c0_n29_w115, 
            w116=> c0_n29_w116, 
            w117=> c0_n29_w117, 
            w118=> c0_n29_w118, 
            w119=> c0_n29_w119, 
            w120=> c0_n29_w120, 
            w121=> c0_n29_w121, 
            w122=> c0_n29_w122, 
            w123=> c0_n29_w123, 
            w124=> c0_n29_w124, 
            w125=> c0_n29_w125, 
            w126=> c0_n29_w126, 
            w127=> c0_n29_w127, 
            w128=> c0_n29_w128, 
            w129=> c0_n29_w129, 
            w130=> c0_n29_w130, 
            w131=> c0_n29_w131, 
            w132=> c0_n29_w132, 
            w133=> c0_n29_w133, 
            w134=> c0_n29_w134, 
            w135=> c0_n29_w135, 
            w136=> c0_n29_w136, 
            w137=> c0_n29_w137, 
            w138=> c0_n29_w138, 
            w139=> c0_n29_w139, 
            w140=> c0_n29_w140, 
            w141=> c0_n29_w141, 
            w142=> c0_n29_w142, 
            w143=> c0_n29_w143, 
            w144=> c0_n29_w144, 
            w145=> c0_n29_w145, 
            w146=> c0_n29_w146, 
            w147=> c0_n29_w147, 
            w148=> c0_n29_w148, 
            w149=> c0_n29_w149, 
            w150=> c0_n29_w150, 
            w151=> c0_n29_w151, 
            w152=> c0_n29_w152, 
            w153=> c0_n29_w153, 
            w154=> c0_n29_w154, 
            w155=> c0_n29_w155, 
            w156=> c0_n29_w156, 
            w157=> c0_n29_w157, 
            w158=> c0_n29_w158, 
            w159=> c0_n29_w159, 
            w160=> c0_n29_w160, 
            w161=> c0_n29_w161, 
            w162=> c0_n29_w162, 
            w163=> c0_n29_w163, 
            w164=> c0_n29_w164, 
            w165=> c0_n29_w165, 
            w166=> c0_n29_w166, 
            w167=> c0_n29_w167, 
            w168=> c0_n29_w168, 
            w169=> c0_n29_w169, 
            w170=> c0_n29_w170, 
            w171=> c0_n29_w171, 
            w172=> c0_n29_w172, 
            w173=> c0_n29_w173, 
            w174=> c0_n29_w174, 
            w175=> c0_n29_w175, 
            w176=> c0_n29_w176, 
            w177=> c0_n29_w177, 
            w178=> c0_n29_w178, 
            w179=> c0_n29_w179, 
            w180=> c0_n29_w180, 
            w181=> c0_n29_w181, 
            w182=> c0_n29_w182, 
            w183=> c0_n29_w183, 
            w184=> c0_n29_w184, 
            w185=> c0_n29_w185, 
            w186=> c0_n29_w186, 
            w187=> c0_n29_w187, 
            w188=> c0_n29_w188, 
            w189=> c0_n29_w189, 
            w190=> c0_n29_w190, 
            w191=> c0_n29_w191, 
            w192=> c0_n29_w192, 
            w193=> c0_n29_w193, 
            w194=> c0_n29_w194, 
            w195=> c0_n29_w195, 
            w196=> c0_n29_w196, 
            w197=> c0_n29_w197, 
            w198=> c0_n29_w198, 
            w199=> c0_n29_w199, 
            w200=> c0_n29_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n29_y
   );           
            
neuron_inst_30: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n30_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n30_w1, 
            w2=> c0_n30_w2, 
            w3=> c0_n30_w3, 
            w4=> c0_n30_w4, 
            w5=> c0_n30_w5, 
            w6=> c0_n30_w6, 
            w7=> c0_n30_w7, 
            w8=> c0_n30_w8, 
            w9=> c0_n30_w9, 
            w10=> c0_n30_w10, 
            w11=> c0_n30_w11, 
            w12=> c0_n30_w12, 
            w13=> c0_n30_w13, 
            w14=> c0_n30_w14, 
            w15=> c0_n30_w15, 
            w16=> c0_n30_w16, 
            w17=> c0_n30_w17, 
            w18=> c0_n30_w18, 
            w19=> c0_n30_w19, 
            w20=> c0_n30_w20, 
            w21=> c0_n30_w21, 
            w22=> c0_n30_w22, 
            w23=> c0_n30_w23, 
            w24=> c0_n30_w24, 
            w25=> c0_n30_w25, 
            w26=> c0_n30_w26, 
            w27=> c0_n30_w27, 
            w28=> c0_n30_w28, 
            w29=> c0_n30_w29, 
            w30=> c0_n30_w30, 
            w31=> c0_n30_w31, 
            w32=> c0_n30_w32, 
            w33=> c0_n30_w33, 
            w34=> c0_n30_w34, 
            w35=> c0_n30_w35, 
            w36=> c0_n30_w36, 
            w37=> c0_n30_w37, 
            w38=> c0_n30_w38, 
            w39=> c0_n30_w39, 
            w40=> c0_n30_w40, 
            w41=> c0_n30_w41, 
            w42=> c0_n30_w42, 
            w43=> c0_n30_w43, 
            w44=> c0_n30_w44, 
            w45=> c0_n30_w45, 
            w46=> c0_n30_w46, 
            w47=> c0_n30_w47, 
            w48=> c0_n30_w48, 
            w49=> c0_n30_w49, 
            w50=> c0_n30_w50, 
            w51=> c0_n30_w51, 
            w52=> c0_n30_w52, 
            w53=> c0_n30_w53, 
            w54=> c0_n30_w54, 
            w55=> c0_n30_w55, 
            w56=> c0_n30_w56, 
            w57=> c0_n30_w57, 
            w58=> c0_n30_w58, 
            w59=> c0_n30_w59, 
            w60=> c0_n30_w60, 
            w61=> c0_n30_w61, 
            w62=> c0_n30_w62, 
            w63=> c0_n30_w63, 
            w64=> c0_n30_w64, 
            w65=> c0_n30_w65, 
            w66=> c0_n30_w66, 
            w67=> c0_n30_w67, 
            w68=> c0_n30_w68, 
            w69=> c0_n30_w69, 
            w70=> c0_n30_w70, 
            w71=> c0_n30_w71, 
            w72=> c0_n30_w72, 
            w73=> c0_n30_w73, 
            w74=> c0_n30_w74, 
            w75=> c0_n30_w75, 
            w76=> c0_n30_w76, 
            w77=> c0_n30_w77, 
            w78=> c0_n30_w78, 
            w79=> c0_n30_w79, 
            w80=> c0_n30_w80, 
            w81=> c0_n30_w81, 
            w82=> c0_n30_w82, 
            w83=> c0_n30_w83, 
            w84=> c0_n30_w84, 
            w85=> c0_n30_w85, 
            w86=> c0_n30_w86, 
            w87=> c0_n30_w87, 
            w88=> c0_n30_w88, 
            w89=> c0_n30_w89, 
            w90=> c0_n30_w90, 
            w91=> c0_n30_w91, 
            w92=> c0_n30_w92, 
            w93=> c0_n30_w93, 
            w94=> c0_n30_w94, 
            w95=> c0_n30_w95, 
            w96=> c0_n30_w96, 
            w97=> c0_n30_w97, 
            w98=> c0_n30_w98, 
            w99=> c0_n30_w99, 
            w100=> c0_n30_w100, 
            w101=> c0_n30_w101, 
            w102=> c0_n30_w102, 
            w103=> c0_n30_w103, 
            w104=> c0_n30_w104, 
            w105=> c0_n30_w105, 
            w106=> c0_n30_w106, 
            w107=> c0_n30_w107, 
            w108=> c0_n30_w108, 
            w109=> c0_n30_w109, 
            w110=> c0_n30_w110, 
            w111=> c0_n30_w111, 
            w112=> c0_n30_w112, 
            w113=> c0_n30_w113, 
            w114=> c0_n30_w114, 
            w115=> c0_n30_w115, 
            w116=> c0_n30_w116, 
            w117=> c0_n30_w117, 
            w118=> c0_n30_w118, 
            w119=> c0_n30_w119, 
            w120=> c0_n30_w120, 
            w121=> c0_n30_w121, 
            w122=> c0_n30_w122, 
            w123=> c0_n30_w123, 
            w124=> c0_n30_w124, 
            w125=> c0_n30_w125, 
            w126=> c0_n30_w126, 
            w127=> c0_n30_w127, 
            w128=> c0_n30_w128, 
            w129=> c0_n30_w129, 
            w130=> c0_n30_w130, 
            w131=> c0_n30_w131, 
            w132=> c0_n30_w132, 
            w133=> c0_n30_w133, 
            w134=> c0_n30_w134, 
            w135=> c0_n30_w135, 
            w136=> c0_n30_w136, 
            w137=> c0_n30_w137, 
            w138=> c0_n30_w138, 
            w139=> c0_n30_w139, 
            w140=> c0_n30_w140, 
            w141=> c0_n30_w141, 
            w142=> c0_n30_w142, 
            w143=> c0_n30_w143, 
            w144=> c0_n30_w144, 
            w145=> c0_n30_w145, 
            w146=> c0_n30_w146, 
            w147=> c0_n30_w147, 
            w148=> c0_n30_w148, 
            w149=> c0_n30_w149, 
            w150=> c0_n30_w150, 
            w151=> c0_n30_w151, 
            w152=> c0_n30_w152, 
            w153=> c0_n30_w153, 
            w154=> c0_n30_w154, 
            w155=> c0_n30_w155, 
            w156=> c0_n30_w156, 
            w157=> c0_n30_w157, 
            w158=> c0_n30_w158, 
            w159=> c0_n30_w159, 
            w160=> c0_n30_w160, 
            w161=> c0_n30_w161, 
            w162=> c0_n30_w162, 
            w163=> c0_n30_w163, 
            w164=> c0_n30_w164, 
            w165=> c0_n30_w165, 
            w166=> c0_n30_w166, 
            w167=> c0_n30_w167, 
            w168=> c0_n30_w168, 
            w169=> c0_n30_w169, 
            w170=> c0_n30_w170, 
            w171=> c0_n30_w171, 
            w172=> c0_n30_w172, 
            w173=> c0_n30_w173, 
            w174=> c0_n30_w174, 
            w175=> c0_n30_w175, 
            w176=> c0_n30_w176, 
            w177=> c0_n30_w177, 
            w178=> c0_n30_w178, 
            w179=> c0_n30_w179, 
            w180=> c0_n30_w180, 
            w181=> c0_n30_w181, 
            w182=> c0_n30_w182, 
            w183=> c0_n30_w183, 
            w184=> c0_n30_w184, 
            w185=> c0_n30_w185, 
            w186=> c0_n30_w186, 
            w187=> c0_n30_w187, 
            w188=> c0_n30_w188, 
            w189=> c0_n30_w189, 
            w190=> c0_n30_w190, 
            w191=> c0_n30_w191, 
            w192=> c0_n30_w192, 
            w193=> c0_n30_w193, 
            w194=> c0_n30_w194, 
            w195=> c0_n30_w195, 
            w196=> c0_n30_w196, 
            w197=> c0_n30_w197, 
            w198=> c0_n30_w198, 
            w199=> c0_n30_w199, 
            w200=> c0_n30_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n30_y
   );           
            
neuron_inst_31: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n31_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n31_w1, 
            w2=> c0_n31_w2, 
            w3=> c0_n31_w3, 
            w4=> c0_n31_w4, 
            w5=> c0_n31_w5, 
            w6=> c0_n31_w6, 
            w7=> c0_n31_w7, 
            w8=> c0_n31_w8, 
            w9=> c0_n31_w9, 
            w10=> c0_n31_w10, 
            w11=> c0_n31_w11, 
            w12=> c0_n31_w12, 
            w13=> c0_n31_w13, 
            w14=> c0_n31_w14, 
            w15=> c0_n31_w15, 
            w16=> c0_n31_w16, 
            w17=> c0_n31_w17, 
            w18=> c0_n31_w18, 
            w19=> c0_n31_w19, 
            w20=> c0_n31_w20, 
            w21=> c0_n31_w21, 
            w22=> c0_n31_w22, 
            w23=> c0_n31_w23, 
            w24=> c0_n31_w24, 
            w25=> c0_n31_w25, 
            w26=> c0_n31_w26, 
            w27=> c0_n31_w27, 
            w28=> c0_n31_w28, 
            w29=> c0_n31_w29, 
            w30=> c0_n31_w30, 
            w31=> c0_n31_w31, 
            w32=> c0_n31_w32, 
            w33=> c0_n31_w33, 
            w34=> c0_n31_w34, 
            w35=> c0_n31_w35, 
            w36=> c0_n31_w36, 
            w37=> c0_n31_w37, 
            w38=> c0_n31_w38, 
            w39=> c0_n31_w39, 
            w40=> c0_n31_w40, 
            w41=> c0_n31_w41, 
            w42=> c0_n31_w42, 
            w43=> c0_n31_w43, 
            w44=> c0_n31_w44, 
            w45=> c0_n31_w45, 
            w46=> c0_n31_w46, 
            w47=> c0_n31_w47, 
            w48=> c0_n31_w48, 
            w49=> c0_n31_w49, 
            w50=> c0_n31_w50, 
            w51=> c0_n31_w51, 
            w52=> c0_n31_w52, 
            w53=> c0_n31_w53, 
            w54=> c0_n31_w54, 
            w55=> c0_n31_w55, 
            w56=> c0_n31_w56, 
            w57=> c0_n31_w57, 
            w58=> c0_n31_w58, 
            w59=> c0_n31_w59, 
            w60=> c0_n31_w60, 
            w61=> c0_n31_w61, 
            w62=> c0_n31_w62, 
            w63=> c0_n31_w63, 
            w64=> c0_n31_w64, 
            w65=> c0_n31_w65, 
            w66=> c0_n31_w66, 
            w67=> c0_n31_w67, 
            w68=> c0_n31_w68, 
            w69=> c0_n31_w69, 
            w70=> c0_n31_w70, 
            w71=> c0_n31_w71, 
            w72=> c0_n31_w72, 
            w73=> c0_n31_w73, 
            w74=> c0_n31_w74, 
            w75=> c0_n31_w75, 
            w76=> c0_n31_w76, 
            w77=> c0_n31_w77, 
            w78=> c0_n31_w78, 
            w79=> c0_n31_w79, 
            w80=> c0_n31_w80, 
            w81=> c0_n31_w81, 
            w82=> c0_n31_w82, 
            w83=> c0_n31_w83, 
            w84=> c0_n31_w84, 
            w85=> c0_n31_w85, 
            w86=> c0_n31_w86, 
            w87=> c0_n31_w87, 
            w88=> c0_n31_w88, 
            w89=> c0_n31_w89, 
            w90=> c0_n31_w90, 
            w91=> c0_n31_w91, 
            w92=> c0_n31_w92, 
            w93=> c0_n31_w93, 
            w94=> c0_n31_w94, 
            w95=> c0_n31_w95, 
            w96=> c0_n31_w96, 
            w97=> c0_n31_w97, 
            w98=> c0_n31_w98, 
            w99=> c0_n31_w99, 
            w100=> c0_n31_w100, 
            w101=> c0_n31_w101, 
            w102=> c0_n31_w102, 
            w103=> c0_n31_w103, 
            w104=> c0_n31_w104, 
            w105=> c0_n31_w105, 
            w106=> c0_n31_w106, 
            w107=> c0_n31_w107, 
            w108=> c0_n31_w108, 
            w109=> c0_n31_w109, 
            w110=> c0_n31_w110, 
            w111=> c0_n31_w111, 
            w112=> c0_n31_w112, 
            w113=> c0_n31_w113, 
            w114=> c0_n31_w114, 
            w115=> c0_n31_w115, 
            w116=> c0_n31_w116, 
            w117=> c0_n31_w117, 
            w118=> c0_n31_w118, 
            w119=> c0_n31_w119, 
            w120=> c0_n31_w120, 
            w121=> c0_n31_w121, 
            w122=> c0_n31_w122, 
            w123=> c0_n31_w123, 
            w124=> c0_n31_w124, 
            w125=> c0_n31_w125, 
            w126=> c0_n31_w126, 
            w127=> c0_n31_w127, 
            w128=> c0_n31_w128, 
            w129=> c0_n31_w129, 
            w130=> c0_n31_w130, 
            w131=> c0_n31_w131, 
            w132=> c0_n31_w132, 
            w133=> c0_n31_w133, 
            w134=> c0_n31_w134, 
            w135=> c0_n31_w135, 
            w136=> c0_n31_w136, 
            w137=> c0_n31_w137, 
            w138=> c0_n31_w138, 
            w139=> c0_n31_w139, 
            w140=> c0_n31_w140, 
            w141=> c0_n31_w141, 
            w142=> c0_n31_w142, 
            w143=> c0_n31_w143, 
            w144=> c0_n31_w144, 
            w145=> c0_n31_w145, 
            w146=> c0_n31_w146, 
            w147=> c0_n31_w147, 
            w148=> c0_n31_w148, 
            w149=> c0_n31_w149, 
            w150=> c0_n31_w150, 
            w151=> c0_n31_w151, 
            w152=> c0_n31_w152, 
            w153=> c0_n31_w153, 
            w154=> c0_n31_w154, 
            w155=> c0_n31_w155, 
            w156=> c0_n31_w156, 
            w157=> c0_n31_w157, 
            w158=> c0_n31_w158, 
            w159=> c0_n31_w159, 
            w160=> c0_n31_w160, 
            w161=> c0_n31_w161, 
            w162=> c0_n31_w162, 
            w163=> c0_n31_w163, 
            w164=> c0_n31_w164, 
            w165=> c0_n31_w165, 
            w166=> c0_n31_w166, 
            w167=> c0_n31_w167, 
            w168=> c0_n31_w168, 
            w169=> c0_n31_w169, 
            w170=> c0_n31_w170, 
            w171=> c0_n31_w171, 
            w172=> c0_n31_w172, 
            w173=> c0_n31_w173, 
            w174=> c0_n31_w174, 
            w175=> c0_n31_w175, 
            w176=> c0_n31_w176, 
            w177=> c0_n31_w177, 
            w178=> c0_n31_w178, 
            w179=> c0_n31_w179, 
            w180=> c0_n31_w180, 
            w181=> c0_n31_w181, 
            w182=> c0_n31_w182, 
            w183=> c0_n31_w183, 
            w184=> c0_n31_w184, 
            w185=> c0_n31_w185, 
            w186=> c0_n31_w186, 
            w187=> c0_n31_w187, 
            w188=> c0_n31_w188, 
            w189=> c0_n31_w189, 
            w190=> c0_n31_w190, 
            w191=> c0_n31_w191, 
            w192=> c0_n31_w192, 
            w193=> c0_n31_w193, 
            w194=> c0_n31_w194, 
            w195=> c0_n31_w195, 
            w196=> c0_n31_w196, 
            w197=> c0_n31_w197, 
            w198=> c0_n31_w198, 
            w199=> c0_n31_w199, 
            w200=> c0_n31_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n31_y
   );           
            
neuron_inst_32: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n32_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n32_w1, 
            w2=> c0_n32_w2, 
            w3=> c0_n32_w3, 
            w4=> c0_n32_w4, 
            w5=> c0_n32_w5, 
            w6=> c0_n32_w6, 
            w7=> c0_n32_w7, 
            w8=> c0_n32_w8, 
            w9=> c0_n32_w9, 
            w10=> c0_n32_w10, 
            w11=> c0_n32_w11, 
            w12=> c0_n32_w12, 
            w13=> c0_n32_w13, 
            w14=> c0_n32_w14, 
            w15=> c0_n32_w15, 
            w16=> c0_n32_w16, 
            w17=> c0_n32_w17, 
            w18=> c0_n32_w18, 
            w19=> c0_n32_w19, 
            w20=> c0_n32_w20, 
            w21=> c0_n32_w21, 
            w22=> c0_n32_w22, 
            w23=> c0_n32_w23, 
            w24=> c0_n32_w24, 
            w25=> c0_n32_w25, 
            w26=> c0_n32_w26, 
            w27=> c0_n32_w27, 
            w28=> c0_n32_w28, 
            w29=> c0_n32_w29, 
            w30=> c0_n32_w30, 
            w31=> c0_n32_w31, 
            w32=> c0_n32_w32, 
            w33=> c0_n32_w33, 
            w34=> c0_n32_w34, 
            w35=> c0_n32_w35, 
            w36=> c0_n32_w36, 
            w37=> c0_n32_w37, 
            w38=> c0_n32_w38, 
            w39=> c0_n32_w39, 
            w40=> c0_n32_w40, 
            w41=> c0_n32_w41, 
            w42=> c0_n32_w42, 
            w43=> c0_n32_w43, 
            w44=> c0_n32_w44, 
            w45=> c0_n32_w45, 
            w46=> c0_n32_w46, 
            w47=> c0_n32_w47, 
            w48=> c0_n32_w48, 
            w49=> c0_n32_w49, 
            w50=> c0_n32_w50, 
            w51=> c0_n32_w51, 
            w52=> c0_n32_w52, 
            w53=> c0_n32_w53, 
            w54=> c0_n32_w54, 
            w55=> c0_n32_w55, 
            w56=> c0_n32_w56, 
            w57=> c0_n32_w57, 
            w58=> c0_n32_w58, 
            w59=> c0_n32_w59, 
            w60=> c0_n32_w60, 
            w61=> c0_n32_w61, 
            w62=> c0_n32_w62, 
            w63=> c0_n32_w63, 
            w64=> c0_n32_w64, 
            w65=> c0_n32_w65, 
            w66=> c0_n32_w66, 
            w67=> c0_n32_w67, 
            w68=> c0_n32_w68, 
            w69=> c0_n32_w69, 
            w70=> c0_n32_w70, 
            w71=> c0_n32_w71, 
            w72=> c0_n32_w72, 
            w73=> c0_n32_w73, 
            w74=> c0_n32_w74, 
            w75=> c0_n32_w75, 
            w76=> c0_n32_w76, 
            w77=> c0_n32_w77, 
            w78=> c0_n32_w78, 
            w79=> c0_n32_w79, 
            w80=> c0_n32_w80, 
            w81=> c0_n32_w81, 
            w82=> c0_n32_w82, 
            w83=> c0_n32_w83, 
            w84=> c0_n32_w84, 
            w85=> c0_n32_w85, 
            w86=> c0_n32_w86, 
            w87=> c0_n32_w87, 
            w88=> c0_n32_w88, 
            w89=> c0_n32_w89, 
            w90=> c0_n32_w90, 
            w91=> c0_n32_w91, 
            w92=> c0_n32_w92, 
            w93=> c0_n32_w93, 
            w94=> c0_n32_w94, 
            w95=> c0_n32_w95, 
            w96=> c0_n32_w96, 
            w97=> c0_n32_w97, 
            w98=> c0_n32_w98, 
            w99=> c0_n32_w99, 
            w100=> c0_n32_w100, 
            w101=> c0_n32_w101, 
            w102=> c0_n32_w102, 
            w103=> c0_n32_w103, 
            w104=> c0_n32_w104, 
            w105=> c0_n32_w105, 
            w106=> c0_n32_w106, 
            w107=> c0_n32_w107, 
            w108=> c0_n32_w108, 
            w109=> c0_n32_w109, 
            w110=> c0_n32_w110, 
            w111=> c0_n32_w111, 
            w112=> c0_n32_w112, 
            w113=> c0_n32_w113, 
            w114=> c0_n32_w114, 
            w115=> c0_n32_w115, 
            w116=> c0_n32_w116, 
            w117=> c0_n32_w117, 
            w118=> c0_n32_w118, 
            w119=> c0_n32_w119, 
            w120=> c0_n32_w120, 
            w121=> c0_n32_w121, 
            w122=> c0_n32_w122, 
            w123=> c0_n32_w123, 
            w124=> c0_n32_w124, 
            w125=> c0_n32_w125, 
            w126=> c0_n32_w126, 
            w127=> c0_n32_w127, 
            w128=> c0_n32_w128, 
            w129=> c0_n32_w129, 
            w130=> c0_n32_w130, 
            w131=> c0_n32_w131, 
            w132=> c0_n32_w132, 
            w133=> c0_n32_w133, 
            w134=> c0_n32_w134, 
            w135=> c0_n32_w135, 
            w136=> c0_n32_w136, 
            w137=> c0_n32_w137, 
            w138=> c0_n32_w138, 
            w139=> c0_n32_w139, 
            w140=> c0_n32_w140, 
            w141=> c0_n32_w141, 
            w142=> c0_n32_w142, 
            w143=> c0_n32_w143, 
            w144=> c0_n32_w144, 
            w145=> c0_n32_w145, 
            w146=> c0_n32_w146, 
            w147=> c0_n32_w147, 
            w148=> c0_n32_w148, 
            w149=> c0_n32_w149, 
            w150=> c0_n32_w150, 
            w151=> c0_n32_w151, 
            w152=> c0_n32_w152, 
            w153=> c0_n32_w153, 
            w154=> c0_n32_w154, 
            w155=> c0_n32_w155, 
            w156=> c0_n32_w156, 
            w157=> c0_n32_w157, 
            w158=> c0_n32_w158, 
            w159=> c0_n32_w159, 
            w160=> c0_n32_w160, 
            w161=> c0_n32_w161, 
            w162=> c0_n32_w162, 
            w163=> c0_n32_w163, 
            w164=> c0_n32_w164, 
            w165=> c0_n32_w165, 
            w166=> c0_n32_w166, 
            w167=> c0_n32_w167, 
            w168=> c0_n32_w168, 
            w169=> c0_n32_w169, 
            w170=> c0_n32_w170, 
            w171=> c0_n32_w171, 
            w172=> c0_n32_w172, 
            w173=> c0_n32_w173, 
            w174=> c0_n32_w174, 
            w175=> c0_n32_w175, 
            w176=> c0_n32_w176, 
            w177=> c0_n32_w177, 
            w178=> c0_n32_w178, 
            w179=> c0_n32_w179, 
            w180=> c0_n32_w180, 
            w181=> c0_n32_w181, 
            w182=> c0_n32_w182, 
            w183=> c0_n32_w183, 
            w184=> c0_n32_w184, 
            w185=> c0_n32_w185, 
            w186=> c0_n32_w186, 
            w187=> c0_n32_w187, 
            w188=> c0_n32_w188, 
            w189=> c0_n32_w189, 
            w190=> c0_n32_w190, 
            w191=> c0_n32_w191, 
            w192=> c0_n32_w192, 
            w193=> c0_n32_w193, 
            w194=> c0_n32_w194, 
            w195=> c0_n32_w195, 
            w196=> c0_n32_w196, 
            w197=> c0_n32_w197, 
            w198=> c0_n32_w198, 
            w199=> c0_n32_w199, 
            w200=> c0_n32_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n32_y
   );           
            
neuron_inst_33: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n33_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n33_w1, 
            w2=> c0_n33_w2, 
            w3=> c0_n33_w3, 
            w4=> c0_n33_w4, 
            w5=> c0_n33_w5, 
            w6=> c0_n33_w6, 
            w7=> c0_n33_w7, 
            w8=> c0_n33_w8, 
            w9=> c0_n33_w9, 
            w10=> c0_n33_w10, 
            w11=> c0_n33_w11, 
            w12=> c0_n33_w12, 
            w13=> c0_n33_w13, 
            w14=> c0_n33_w14, 
            w15=> c0_n33_w15, 
            w16=> c0_n33_w16, 
            w17=> c0_n33_w17, 
            w18=> c0_n33_w18, 
            w19=> c0_n33_w19, 
            w20=> c0_n33_w20, 
            w21=> c0_n33_w21, 
            w22=> c0_n33_w22, 
            w23=> c0_n33_w23, 
            w24=> c0_n33_w24, 
            w25=> c0_n33_w25, 
            w26=> c0_n33_w26, 
            w27=> c0_n33_w27, 
            w28=> c0_n33_w28, 
            w29=> c0_n33_w29, 
            w30=> c0_n33_w30, 
            w31=> c0_n33_w31, 
            w32=> c0_n33_w32, 
            w33=> c0_n33_w33, 
            w34=> c0_n33_w34, 
            w35=> c0_n33_w35, 
            w36=> c0_n33_w36, 
            w37=> c0_n33_w37, 
            w38=> c0_n33_w38, 
            w39=> c0_n33_w39, 
            w40=> c0_n33_w40, 
            w41=> c0_n33_w41, 
            w42=> c0_n33_w42, 
            w43=> c0_n33_w43, 
            w44=> c0_n33_w44, 
            w45=> c0_n33_w45, 
            w46=> c0_n33_w46, 
            w47=> c0_n33_w47, 
            w48=> c0_n33_w48, 
            w49=> c0_n33_w49, 
            w50=> c0_n33_w50, 
            w51=> c0_n33_w51, 
            w52=> c0_n33_w52, 
            w53=> c0_n33_w53, 
            w54=> c0_n33_w54, 
            w55=> c0_n33_w55, 
            w56=> c0_n33_w56, 
            w57=> c0_n33_w57, 
            w58=> c0_n33_w58, 
            w59=> c0_n33_w59, 
            w60=> c0_n33_w60, 
            w61=> c0_n33_w61, 
            w62=> c0_n33_w62, 
            w63=> c0_n33_w63, 
            w64=> c0_n33_w64, 
            w65=> c0_n33_w65, 
            w66=> c0_n33_w66, 
            w67=> c0_n33_w67, 
            w68=> c0_n33_w68, 
            w69=> c0_n33_w69, 
            w70=> c0_n33_w70, 
            w71=> c0_n33_w71, 
            w72=> c0_n33_w72, 
            w73=> c0_n33_w73, 
            w74=> c0_n33_w74, 
            w75=> c0_n33_w75, 
            w76=> c0_n33_w76, 
            w77=> c0_n33_w77, 
            w78=> c0_n33_w78, 
            w79=> c0_n33_w79, 
            w80=> c0_n33_w80, 
            w81=> c0_n33_w81, 
            w82=> c0_n33_w82, 
            w83=> c0_n33_w83, 
            w84=> c0_n33_w84, 
            w85=> c0_n33_w85, 
            w86=> c0_n33_w86, 
            w87=> c0_n33_w87, 
            w88=> c0_n33_w88, 
            w89=> c0_n33_w89, 
            w90=> c0_n33_w90, 
            w91=> c0_n33_w91, 
            w92=> c0_n33_w92, 
            w93=> c0_n33_w93, 
            w94=> c0_n33_w94, 
            w95=> c0_n33_w95, 
            w96=> c0_n33_w96, 
            w97=> c0_n33_w97, 
            w98=> c0_n33_w98, 
            w99=> c0_n33_w99, 
            w100=> c0_n33_w100, 
            w101=> c0_n33_w101, 
            w102=> c0_n33_w102, 
            w103=> c0_n33_w103, 
            w104=> c0_n33_w104, 
            w105=> c0_n33_w105, 
            w106=> c0_n33_w106, 
            w107=> c0_n33_w107, 
            w108=> c0_n33_w108, 
            w109=> c0_n33_w109, 
            w110=> c0_n33_w110, 
            w111=> c0_n33_w111, 
            w112=> c0_n33_w112, 
            w113=> c0_n33_w113, 
            w114=> c0_n33_w114, 
            w115=> c0_n33_w115, 
            w116=> c0_n33_w116, 
            w117=> c0_n33_w117, 
            w118=> c0_n33_w118, 
            w119=> c0_n33_w119, 
            w120=> c0_n33_w120, 
            w121=> c0_n33_w121, 
            w122=> c0_n33_w122, 
            w123=> c0_n33_w123, 
            w124=> c0_n33_w124, 
            w125=> c0_n33_w125, 
            w126=> c0_n33_w126, 
            w127=> c0_n33_w127, 
            w128=> c0_n33_w128, 
            w129=> c0_n33_w129, 
            w130=> c0_n33_w130, 
            w131=> c0_n33_w131, 
            w132=> c0_n33_w132, 
            w133=> c0_n33_w133, 
            w134=> c0_n33_w134, 
            w135=> c0_n33_w135, 
            w136=> c0_n33_w136, 
            w137=> c0_n33_w137, 
            w138=> c0_n33_w138, 
            w139=> c0_n33_w139, 
            w140=> c0_n33_w140, 
            w141=> c0_n33_w141, 
            w142=> c0_n33_w142, 
            w143=> c0_n33_w143, 
            w144=> c0_n33_w144, 
            w145=> c0_n33_w145, 
            w146=> c0_n33_w146, 
            w147=> c0_n33_w147, 
            w148=> c0_n33_w148, 
            w149=> c0_n33_w149, 
            w150=> c0_n33_w150, 
            w151=> c0_n33_w151, 
            w152=> c0_n33_w152, 
            w153=> c0_n33_w153, 
            w154=> c0_n33_w154, 
            w155=> c0_n33_w155, 
            w156=> c0_n33_w156, 
            w157=> c0_n33_w157, 
            w158=> c0_n33_w158, 
            w159=> c0_n33_w159, 
            w160=> c0_n33_w160, 
            w161=> c0_n33_w161, 
            w162=> c0_n33_w162, 
            w163=> c0_n33_w163, 
            w164=> c0_n33_w164, 
            w165=> c0_n33_w165, 
            w166=> c0_n33_w166, 
            w167=> c0_n33_w167, 
            w168=> c0_n33_w168, 
            w169=> c0_n33_w169, 
            w170=> c0_n33_w170, 
            w171=> c0_n33_w171, 
            w172=> c0_n33_w172, 
            w173=> c0_n33_w173, 
            w174=> c0_n33_w174, 
            w175=> c0_n33_w175, 
            w176=> c0_n33_w176, 
            w177=> c0_n33_w177, 
            w178=> c0_n33_w178, 
            w179=> c0_n33_w179, 
            w180=> c0_n33_w180, 
            w181=> c0_n33_w181, 
            w182=> c0_n33_w182, 
            w183=> c0_n33_w183, 
            w184=> c0_n33_w184, 
            w185=> c0_n33_w185, 
            w186=> c0_n33_w186, 
            w187=> c0_n33_w187, 
            w188=> c0_n33_w188, 
            w189=> c0_n33_w189, 
            w190=> c0_n33_w190, 
            w191=> c0_n33_w191, 
            w192=> c0_n33_w192, 
            w193=> c0_n33_w193, 
            w194=> c0_n33_w194, 
            w195=> c0_n33_w195, 
            w196=> c0_n33_w196, 
            w197=> c0_n33_w197, 
            w198=> c0_n33_w198, 
            w199=> c0_n33_w199, 
            w200=> c0_n33_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n33_y
   );           
            
neuron_inst_34: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n34_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n34_w1, 
            w2=> c0_n34_w2, 
            w3=> c0_n34_w3, 
            w4=> c0_n34_w4, 
            w5=> c0_n34_w5, 
            w6=> c0_n34_w6, 
            w7=> c0_n34_w7, 
            w8=> c0_n34_w8, 
            w9=> c0_n34_w9, 
            w10=> c0_n34_w10, 
            w11=> c0_n34_w11, 
            w12=> c0_n34_w12, 
            w13=> c0_n34_w13, 
            w14=> c0_n34_w14, 
            w15=> c0_n34_w15, 
            w16=> c0_n34_w16, 
            w17=> c0_n34_w17, 
            w18=> c0_n34_w18, 
            w19=> c0_n34_w19, 
            w20=> c0_n34_w20, 
            w21=> c0_n34_w21, 
            w22=> c0_n34_w22, 
            w23=> c0_n34_w23, 
            w24=> c0_n34_w24, 
            w25=> c0_n34_w25, 
            w26=> c0_n34_w26, 
            w27=> c0_n34_w27, 
            w28=> c0_n34_w28, 
            w29=> c0_n34_w29, 
            w30=> c0_n34_w30, 
            w31=> c0_n34_w31, 
            w32=> c0_n34_w32, 
            w33=> c0_n34_w33, 
            w34=> c0_n34_w34, 
            w35=> c0_n34_w35, 
            w36=> c0_n34_w36, 
            w37=> c0_n34_w37, 
            w38=> c0_n34_w38, 
            w39=> c0_n34_w39, 
            w40=> c0_n34_w40, 
            w41=> c0_n34_w41, 
            w42=> c0_n34_w42, 
            w43=> c0_n34_w43, 
            w44=> c0_n34_w44, 
            w45=> c0_n34_w45, 
            w46=> c0_n34_w46, 
            w47=> c0_n34_w47, 
            w48=> c0_n34_w48, 
            w49=> c0_n34_w49, 
            w50=> c0_n34_w50, 
            w51=> c0_n34_w51, 
            w52=> c0_n34_w52, 
            w53=> c0_n34_w53, 
            w54=> c0_n34_w54, 
            w55=> c0_n34_w55, 
            w56=> c0_n34_w56, 
            w57=> c0_n34_w57, 
            w58=> c0_n34_w58, 
            w59=> c0_n34_w59, 
            w60=> c0_n34_w60, 
            w61=> c0_n34_w61, 
            w62=> c0_n34_w62, 
            w63=> c0_n34_w63, 
            w64=> c0_n34_w64, 
            w65=> c0_n34_w65, 
            w66=> c0_n34_w66, 
            w67=> c0_n34_w67, 
            w68=> c0_n34_w68, 
            w69=> c0_n34_w69, 
            w70=> c0_n34_w70, 
            w71=> c0_n34_w71, 
            w72=> c0_n34_w72, 
            w73=> c0_n34_w73, 
            w74=> c0_n34_w74, 
            w75=> c0_n34_w75, 
            w76=> c0_n34_w76, 
            w77=> c0_n34_w77, 
            w78=> c0_n34_w78, 
            w79=> c0_n34_w79, 
            w80=> c0_n34_w80, 
            w81=> c0_n34_w81, 
            w82=> c0_n34_w82, 
            w83=> c0_n34_w83, 
            w84=> c0_n34_w84, 
            w85=> c0_n34_w85, 
            w86=> c0_n34_w86, 
            w87=> c0_n34_w87, 
            w88=> c0_n34_w88, 
            w89=> c0_n34_w89, 
            w90=> c0_n34_w90, 
            w91=> c0_n34_w91, 
            w92=> c0_n34_w92, 
            w93=> c0_n34_w93, 
            w94=> c0_n34_w94, 
            w95=> c0_n34_w95, 
            w96=> c0_n34_w96, 
            w97=> c0_n34_w97, 
            w98=> c0_n34_w98, 
            w99=> c0_n34_w99, 
            w100=> c0_n34_w100, 
            w101=> c0_n34_w101, 
            w102=> c0_n34_w102, 
            w103=> c0_n34_w103, 
            w104=> c0_n34_w104, 
            w105=> c0_n34_w105, 
            w106=> c0_n34_w106, 
            w107=> c0_n34_w107, 
            w108=> c0_n34_w108, 
            w109=> c0_n34_w109, 
            w110=> c0_n34_w110, 
            w111=> c0_n34_w111, 
            w112=> c0_n34_w112, 
            w113=> c0_n34_w113, 
            w114=> c0_n34_w114, 
            w115=> c0_n34_w115, 
            w116=> c0_n34_w116, 
            w117=> c0_n34_w117, 
            w118=> c0_n34_w118, 
            w119=> c0_n34_w119, 
            w120=> c0_n34_w120, 
            w121=> c0_n34_w121, 
            w122=> c0_n34_w122, 
            w123=> c0_n34_w123, 
            w124=> c0_n34_w124, 
            w125=> c0_n34_w125, 
            w126=> c0_n34_w126, 
            w127=> c0_n34_w127, 
            w128=> c0_n34_w128, 
            w129=> c0_n34_w129, 
            w130=> c0_n34_w130, 
            w131=> c0_n34_w131, 
            w132=> c0_n34_w132, 
            w133=> c0_n34_w133, 
            w134=> c0_n34_w134, 
            w135=> c0_n34_w135, 
            w136=> c0_n34_w136, 
            w137=> c0_n34_w137, 
            w138=> c0_n34_w138, 
            w139=> c0_n34_w139, 
            w140=> c0_n34_w140, 
            w141=> c0_n34_w141, 
            w142=> c0_n34_w142, 
            w143=> c0_n34_w143, 
            w144=> c0_n34_w144, 
            w145=> c0_n34_w145, 
            w146=> c0_n34_w146, 
            w147=> c0_n34_w147, 
            w148=> c0_n34_w148, 
            w149=> c0_n34_w149, 
            w150=> c0_n34_w150, 
            w151=> c0_n34_w151, 
            w152=> c0_n34_w152, 
            w153=> c0_n34_w153, 
            w154=> c0_n34_w154, 
            w155=> c0_n34_w155, 
            w156=> c0_n34_w156, 
            w157=> c0_n34_w157, 
            w158=> c0_n34_w158, 
            w159=> c0_n34_w159, 
            w160=> c0_n34_w160, 
            w161=> c0_n34_w161, 
            w162=> c0_n34_w162, 
            w163=> c0_n34_w163, 
            w164=> c0_n34_w164, 
            w165=> c0_n34_w165, 
            w166=> c0_n34_w166, 
            w167=> c0_n34_w167, 
            w168=> c0_n34_w168, 
            w169=> c0_n34_w169, 
            w170=> c0_n34_w170, 
            w171=> c0_n34_w171, 
            w172=> c0_n34_w172, 
            w173=> c0_n34_w173, 
            w174=> c0_n34_w174, 
            w175=> c0_n34_w175, 
            w176=> c0_n34_w176, 
            w177=> c0_n34_w177, 
            w178=> c0_n34_w178, 
            w179=> c0_n34_w179, 
            w180=> c0_n34_w180, 
            w181=> c0_n34_w181, 
            w182=> c0_n34_w182, 
            w183=> c0_n34_w183, 
            w184=> c0_n34_w184, 
            w185=> c0_n34_w185, 
            w186=> c0_n34_w186, 
            w187=> c0_n34_w187, 
            w188=> c0_n34_w188, 
            w189=> c0_n34_w189, 
            w190=> c0_n34_w190, 
            w191=> c0_n34_w191, 
            w192=> c0_n34_w192, 
            w193=> c0_n34_w193, 
            w194=> c0_n34_w194, 
            w195=> c0_n34_w195, 
            w196=> c0_n34_w196, 
            w197=> c0_n34_w197, 
            w198=> c0_n34_w198, 
            w199=> c0_n34_w199, 
            w200=> c0_n34_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n34_y
   );           
            
neuron_inst_35: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n35_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n35_w1, 
            w2=> c0_n35_w2, 
            w3=> c0_n35_w3, 
            w4=> c0_n35_w4, 
            w5=> c0_n35_w5, 
            w6=> c0_n35_w6, 
            w7=> c0_n35_w7, 
            w8=> c0_n35_w8, 
            w9=> c0_n35_w9, 
            w10=> c0_n35_w10, 
            w11=> c0_n35_w11, 
            w12=> c0_n35_w12, 
            w13=> c0_n35_w13, 
            w14=> c0_n35_w14, 
            w15=> c0_n35_w15, 
            w16=> c0_n35_w16, 
            w17=> c0_n35_w17, 
            w18=> c0_n35_w18, 
            w19=> c0_n35_w19, 
            w20=> c0_n35_w20, 
            w21=> c0_n35_w21, 
            w22=> c0_n35_w22, 
            w23=> c0_n35_w23, 
            w24=> c0_n35_w24, 
            w25=> c0_n35_w25, 
            w26=> c0_n35_w26, 
            w27=> c0_n35_w27, 
            w28=> c0_n35_w28, 
            w29=> c0_n35_w29, 
            w30=> c0_n35_w30, 
            w31=> c0_n35_w31, 
            w32=> c0_n35_w32, 
            w33=> c0_n35_w33, 
            w34=> c0_n35_w34, 
            w35=> c0_n35_w35, 
            w36=> c0_n35_w36, 
            w37=> c0_n35_w37, 
            w38=> c0_n35_w38, 
            w39=> c0_n35_w39, 
            w40=> c0_n35_w40, 
            w41=> c0_n35_w41, 
            w42=> c0_n35_w42, 
            w43=> c0_n35_w43, 
            w44=> c0_n35_w44, 
            w45=> c0_n35_w45, 
            w46=> c0_n35_w46, 
            w47=> c0_n35_w47, 
            w48=> c0_n35_w48, 
            w49=> c0_n35_w49, 
            w50=> c0_n35_w50, 
            w51=> c0_n35_w51, 
            w52=> c0_n35_w52, 
            w53=> c0_n35_w53, 
            w54=> c0_n35_w54, 
            w55=> c0_n35_w55, 
            w56=> c0_n35_w56, 
            w57=> c0_n35_w57, 
            w58=> c0_n35_w58, 
            w59=> c0_n35_w59, 
            w60=> c0_n35_w60, 
            w61=> c0_n35_w61, 
            w62=> c0_n35_w62, 
            w63=> c0_n35_w63, 
            w64=> c0_n35_w64, 
            w65=> c0_n35_w65, 
            w66=> c0_n35_w66, 
            w67=> c0_n35_w67, 
            w68=> c0_n35_w68, 
            w69=> c0_n35_w69, 
            w70=> c0_n35_w70, 
            w71=> c0_n35_w71, 
            w72=> c0_n35_w72, 
            w73=> c0_n35_w73, 
            w74=> c0_n35_w74, 
            w75=> c0_n35_w75, 
            w76=> c0_n35_w76, 
            w77=> c0_n35_w77, 
            w78=> c0_n35_w78, 
            w79=> c0_n35_w79, 
            w80=> c0_n35_w80, 
            w81=> c0_n35_w81, 
            w82=> c0_n35_w82, 
            w83=> c0_n35_w83, 
            w84=> c0_n35_w84, 
            w85=> c0_n35_w85, 
            w86=> c0_n35_w86, 
            w87=> c0_n35_w87, 
            w88=> c0_n35_w88, 
            w89=> c0_n35_w89, 
            w90=> c0_n35_w90, 
            w91=> c0_n35_w91, 
            w92=> c0_n35_w92, 
            w93=> c0_n35_w93, 
            w94=> c0_n35_w94, 
            w95=> c0_n35_w95, 
            w96=> c0_n35_w96, 
            w97=> c0_n35_w97, 
            w98=> c0_n35_w98, 
            w99=> c0_n35_w99, 
            w100=> c0_n35_w100, 
            w101=> c0_n35_w101, 
            w102=> c0_n35_w102, 
            w103=> c0_n35_w103, 
            w104=> c0_n35_w104, 
            w105=> c0_n35_w105, 
            w106=> c0_n35_w106, 
            w107=> c0_n35_w107, 
            w108=> c0_n35_w108, 
            w109=> c0_n35_w109, 
            w110=> c0_n35_w110, 
            w111=> c0_n35_w111, 
            w112=> c0_n35_w112, 
            w113=> c0_n35_w113, 
            w114=> c0_n35_w114, 
            w115=> c0_n35_w115, 
            w116=> c0_n35_w116, 
            w117=> c0_n35_w117, 
            w118=> c0_n35_w118, 
            w119=> c0_n35_w119, 
            w120=> c0_n35_w120, 
            w121=> c0_n35_w121, 
            w122=> c0_n35_w122, 
            w123=> c0_n35_w123, 
            w124=> c0_n35_w124, 
            w125=> c0_n35_w125, 
            w126=> c0_n35_w126, 
            w127=> c0_n35_w127, 
            w128=> c0_n35_w128, 
            w129=> c0_n35_w129, 
            w130=> c0_n35_w130, 
            w131=> c0_n35_w131, 
            w132=> c0_n35_w132, 
            w133=> c0_n35_w133, 
            w134=> c0_n35_w134, 
            w135=> c0_n35_w135, 
            w136=> c0_n35_w136, 
            w137=> c0_n35_w137, 
            w138=> c0_n35_w138, 
            w139=> c0_n35_w139, 
            w140=> c0_n35_w140, 
            w141=> c0_n35_w141, 
            w142=> c0_n35_w142, 
            w143=> c0_n35_w143, 
            w144=> c0_n35_w144, 
            w145=> c0_n35_w145, 
            w146=> c0_n35_w146, 
            w147=> c0_n35_w147, 
            w148=> c0_n35_w148, 
            w149=> c0_n35_w149, 
            w150=> c0_n35_w150, 
            w151=> c0_n35_w151, 
            w152=> c0_n35_w152, 
            w153=> c0_n35_w153, 
            w154=> c0_n35_w154, 
            w155=> c0_n35_w155, 
            w156=> c0_n35_w156, 
            w157=> c0_n35_w157, 
            w158=> c0_n35_w158, 
            w159=> c0_n35_w159, 
            w160=> c0_n35_w160, 
            w161=> c0_n35_w161, 
            w162=> c0_n35_w162, 
            w163=> c0_n35_w163, 
            w164=> c0_n35_w164, 
            w165=> c0_n35_w165, 
            w166=> c0_n35_w166, 
            w167=> c0_n35_w167, 
            w168=> c0_n35_w168, 
            w169=> c0_n35_w169, 
            w170=> c0_n35_w170, 
            w171=> c0_n35_w171, 
            w172=> c0_n35_w172, 
            w173=> c0_n35_w173, 
            w174=> c0_n35_w174, 
            w175=> c0_n35_w175, 
            w176=> c0_n35_w176, 
            w177=> c0_n35_w177, 
            w178=> c0_n35_w178, 
            w179=> c0_n35_w179, 
            w180=> c0_n35_w180, 
            w181=> c0_n35_w181, 
            w182=> c0_n35_w182, 
            w183=> c0_n35_w183, 
            w184=> c0_n35_w184, 
            w185=> c0_n35_w185, 
            w186=> c0_n35_w186, 
            w187=> c0_n35_w187, 
            w188=> c0_n35_w188, 
            w189=> c0_n35_w189, 
            w190=> c0_n35_w190, 
            w191=> c0_n35_w191, 
            w192=> c0_n35_w192, 
            w193=> c0_n35_w193, 
            w194=> c0_n35_w194, 
            w195=> c0_n35_w195, 
            w196=> c0_n35_w196, 
            w197=> c0_n35_w197, 
            w198=> c0_n35_w198, 
            w199=> c0_n35_w199, 
            w200=> c0_n35_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n35_y
   );           
            
neuron_inst_36: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n36_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n36_w1, 
            w2=> c0_n36_w2, 
            w3=> c0_n36_w3, 
            w4=> c0_n36_w4, 
            w5=> c0_n36_w5, 
            w6=> c0_n36_w6, 
            w7=> c0_n36_w7, 
            w8=> c0_n36_w8, 
            w9=> c0_n36_w9, 
            w10=> c0_n36_w10, 
            w11=> c0_n36_w11, 
            w12=> c0_n36_w12, 
            w13=> c0_n36_w13, 
            w14=> c0_n36_w14, 
            w15=> c0_n36_w15, 
            w16=> c0_n36_w16, 
            w17=> c0_n36_w17, 
            w18=> c0_n36_w18, 
            w19=> c0_n36_w19, 
            w20=> c0_n36_w20, 
            w21=> c0_n36_w21, 
            w22=> c0_n36_w22, 
            w23=> c0_n36_w23, 
            w24=> c0_n36_w24, 
            w25=> c0_n36_w25, 
            w26=> c0_n36_w26, 
            w27=> c0_n36_w27, 
            w28=> c0_n36_w28, 
            w29=> c0_n36_w29, 
            w30=> c0_n36_w30, 
            w31=> c0_n36_w31, 
            w32=> c0_n36_w32, 
            w33=> c0_n36_w33, 
            w34=> c0_n36_w34, 
            w35=> c0_n36_w35, 
            w36=> c0_n36_w36, 
            w37=> c0_n36_w37, 
            w38=> c0_n36_w38, 
            w39=> c0_n36_w39, 
            w40=> c0_n36_w40, 
            w41=> c0_n36_w41, 
            w42=> c0_n36_w42, 
            w43=> c0_n36_w43, 
            w44=> c0_n36_w44, 
            w45=> c0_n36_w45, 
            w46=> c0_n36_w46, 
            w47=> c0_n36_w47, 
            w48=> c0_n36_w48, 
            w49=> c0_n36_w49, 
            w50=> c0_n36_w50, 
            w51=> c0_n36_w51, 
            w52=> c0_n36_w52, 
            w53=> c0_n36_w53, 
            w54=> c0_n36_w54, 
            w55=> c0_n36_w55, 
            w56=> c0_n36_w56, 
            w57=> c0_n36_w57, 
            w58=> c0_n36_w58, 
            w59=> c0_n36_w59, 
            w60=> c0_n36_w60, 
            w61=> c0_n36_w61, 
            w62=> c0_n36_w62, 
            w63=> c0_n36_w63, 
            w64=> c0_n36_w64, 
            w65=> c0_n36_w65, 
            w66=> c0_n36_w66, 
            w67=> c0_n36_w67, 
            w68=> c0_n36_w68, 
            w69=> c0_n36_w69, 
            w70=> c0_n36_w70, 
            w71=> c0_n36_w71, 
            w72=> c0_n36_w72, 
            w73=> c0_n36_w73, 
            w74=> c0_n36_w74, 
            w75=> c0_n36_w75, 
            w76=> c0_n36_w76, 
            w77=> c0_n36_w77, 
            w78=> c0_n36_w78, 
            w79=> c0_n36_w79, 
            w80=> c0_n36_w80, 
            w81=> c0_n36_w81, 
            w82=> c0_n36_w82, 
            w83=> c0_n36_w83, 
            w84=> c0_n36_w84, 
            w85=> c0_n36_w85, 
            w86=> c0_n36_w86, 
            w87=> c0_n36_w87, 
            w88=> c0_n36_w88, 
            w89=> c0_n36_w89, 
            w90=> c0_n36_w90, 
            w91=> c0_n36_w91, 
            w92=> c0_n36_w92, 
            w93=> c0_n36_w93, 
            w94=> c0_n36_w94, 
            w95=> c0_n36_w95, 
            w96=> c0_n36_w96, 
            w97=> c0_n36_w97, 
            w98=> c0_n36_w98, 
            w99=> c0_n36_w99, 
            w100=> c0_n36_w100, 
            w101=> c0_n36_w101, 
            w102=> c0_n36_w102, 
            w103=> c0_n36_w103, 
            w104=> c0_n36_w104, 
            w105=> c0_n36_w105, 
            w106=> c0_n36_w106, 
            w107=> c0_n36_w107, 
            w108=> c0_n36_w108, 
            w109=> c0_n36_w109, 
            w110=> c0_n36_w110, 
            w111=> c0_n36_w111, 
            w112=> c0_n36_w112, 
            w113=> c0_n36_w113, 
            w114=> c0_n36_w114, 
            w115=> c0_n36_w115, 
            w116=> c0_n36_w116, 
            w117=> c0_n36_w117, 
            w118=> c0_n36_w118, 
            w119=> c0_n36_w119, 
            w120=> c0_n36_w120, 
            w121=> c0_n36_w121, 
            w122=> c0_n36_w122, 
            w123=> c0_n36_w123, 
            w124=> c0_n36_w124, 
            w125=> c0_n36_w125, 
            w126=> c0_n36_w126, 
            w127=> c0_n36_w127, 
            w128=> c0_n36_w128, 
            w129=> c0_n36_w129, 
            w130=> c0_n36_w130, 
            w131=> c0_n36_w131, 
            w132=> c0_n36_w132, 
            w133=> c0_n36_w133, 
            w134=> c0_n36_w134, 
            w135=> c0_n36_w135, 
            w136=> c0_n36_w136, 
            w137=> c0_n36_w137, 
            w138=> c0_n36_w138, 
            w139=> c0_n36_w139, 
            w140=> c0_n36_w140, 
            w141=> c0_n36_w141, 
            w142=> c0_n36_w142, 
            w143=> c0_n36_w143, 
            w144=> c0_n36_w144, 
            w145=> c0_n36_w145, 
            w146=> c0_n36_w146, 
            w147=> c0_n36_w147, 
            w148=> c0_n36_w148, 
            w149=> c0_n36_w149, 
            w150=> c0_n36_w150, 
            w151=> c0_n36_w151, 
            w152=> c0_n36_w152, 
            w153=> c0_n36_w153, 
            w154=> c0_n36_w154, 
            w155=> c0_n36_w155, 
            w156=> c0_n36_w156, 
            w157=> c0_n36_w157, 
            w158=> c0_n36_w158, 
            w159=> c0_n36_w159, 
            w160=> c0_n36_w160, 
            w161=> c0_n36_w161, 
            w162=> c0_n36_w162, 
            w163=> c0_n36_w163, 
            w164=> c0_n36_w164, 
            w165=> c0_n36_w165, 
            w166=> c0_n36_w166, 
            w167=> c0_n36_w167, 
            w168=> c0_n36_w168, 
            w169=> c0_n36_w169, 
            w170=> c0_n36_w170, 
            w171=> c0_n36_w171, 
            w172=> c0_n36_w172, 
            w173=> c0_n36_w173, 
            w174=> c0_n36_w174, 
            w175=> c0_n36_w175, 
            w176=> c0_n36_w176, 
            w177=> c0_n36_w177, 
            w178=> c0_n36_w178, 
            w179=> c0_n36_w179, 
            w180=> c0_n36_w180, 
            w181=> c0_n36_w181, 
            w182=> c0_n36_w182, 
            w183=> c0_n36_w183, 
            w184=> c0_n36_w184, 
            w185=> c0_n36_w185, 
            w186=> c0_n36_w186, 
            w187=> c0_n36_w187, 
            w188=> c0_n36_w188, 
            w189=> c0_n36_w189, 
            w190=> c0_n36_w190, 
            w191=> c0_n36_w191, 
            w192=> c0_n36_w192, 
            w193=> c0_n36_w193, 
            w194=> c0_n36_w194, 
            w195=> c0_n36_w195, 
            w196=> c0_n36_w196, 
            w197=> c0_n36_w197, 
            w198=> c0_n36_w198, 
            w199=> c0_n36_w199, 
            w200=> c0_n36_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n36_y
   );           
            
neuron_inst_37: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n37_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n37_w1, 
            w2=> c0_n37_w2, 
            w3=> c0_n37_w3, 
            w4=> c0_n37_w4, 
            w5=> c0_n37_w5, 
            w6=> c0_n37_w6, 
            w7=> c0_n37_w7, 
            w8=> c0_n37_w8, 
            w9=> c0_n37_w9, 
            w10=> c0_n37_w10, 
            w11=> c0_n37_w11, 
            w12=> c0_n37_w12, 
            w13=> c0_n37_w13, 
            w14=> c0_n37_w14, 
            w15=> c0_n37_w15, 
            w16=> c0_n37_w16, 
            w17=> c0_n37_w17, 
            w18=> c0_n37_w18, 
            w19=> c0_n37_w19, 
            w20=> c0_n37_w20, 
            w21=> c0_n37_w21, 
            w22=> c0_n37_w22, 
            w23=> c0_n37_w23, 
            w24=> c0_n37_w24, 
            w25=> c0_n37_w25, 
            w26=> c0_n37_w26, 
            w27=> c0_n37_w27, 
            w28=> c0_n37_w28, 
            w29=> c0_n37_w29, 
            w30=> c0_n37_w30, 
            w31=> c0_n37_w31, 
            w32=> c0_n37_w32, 
            w33=> c0_n37_w33, 
            w34=> c0_n37_w34, 
            w35=> c0_n37_w35, 
            w36=> c0_n37_w36, 
            w37=> c0_n37_w37, 
            w38=> c0_n37_w38, 
            w39=> c0_n37_w39, 
            w40=> c0_n37_w40, 
            w41=> c0_n37_w41, 
            w42=> c0_n37_w42, 
            w43=> c0_n37_w43, 
            w44=> c0_n37_w44, 
            w45=> c0_n37_w45, 
            w46=> c0_n37_w46, 
            w47=> c0_n37_w47, 
            w48=> c0_n37_w48, 
            w49=> c0_n37_w49, 
            w50=> c0_n37_w50, 
            w51=> c0_n37_w51, 
            w52=> c0_n37_w52, 
            w53=> c0_n37_w53, 
            w54=> c0_n37_w54, 
            w55=> c0_n37_w55, 
            w56=> c0_n37_w56, 
            w57=> c0_n37_w57, 
            w58=> c0_n37_w58, 
            w59=> c0_n37_w59, 
            w60=> c0_n37_w60, 
            w61=> c0_n37_w61, 
            w62=> c0_n37_w62, 
            w63=> c0_n37_w63, 
            w64=> c0_n37_w64, 
            w65=> c0_n37_w65, 
            w66=> c0_n37_w66, 
            w67=> c0_n37_w67, 
            w68=> c0_n37_w68, 
            w69=> c0_n37_w69, 
            w70=> c0_n37_w70, 
            w71=> c0_n37_w71, 
            w72=> c0_n37_w72, 
            w73=> c0_n37_w73, 
            w74=> c0_n37_w74, 
            w75=> c0_n37_w75, 
            w76=> c0_n37_w76, 
            w77=> c0_n37_w77, 
            w78=> c0_n37_w78, 
            w79=> c0_n37_w79, 
            w80=> c0_n37_w80, 
            w81=> c0_n37_w81, 
            w82=> c0_n37_w82, 
            w83=> c0_n37_w83, 
            w84=> c0_n37_w84, 
            w85=> c0_n37_w85, 
            w86=> c0_n37_w86, 
            w87=> c0_n37_w87, 
            w88=> c0_n37_w88, 
            w89=> c0_n37_w89, 
            w90=> c0_n37_w90, 
            w91=> c0_n37_w91, 
            w92=> c0_n37_w92, 
            w93=> c0_n37_w93, 
            w94=> c0_n37_w94, 
            w95=> c0_n37_w95, 
            w96=> c0_n37_w96, 
            w97=> c0_n37_w97, 
            w98=> c0_n37_w98, 
            w99=> c0_n37_w99, 
            w100=> c0_n37_w100, 
            w101=> c0_n37_w101, 
            w102=> c0_n37_w102, 
            w103=> c0_n37_w103, 
            w104=> c0_n37_w104, 
            w105=> c0_n37_w105, 
            w106=> c0_n37_w106, 
            w107=> c0_n37_w107, 
            w108=> c0_n37_w108, 
            w109=> c0_n37_w109, 
            w110=> c0_n37_w110, 
            w111=> c0_n37_w111, 
            w112=> c0_n37_w112, 
            w113=> c0_n37_w113, 
            w114=> c0_n37_w114, 
            w115=> c0_n37_w115, 
            w116=> c0_n37_w116, 
            w117=> c0_n37_w117, 
            w118=> c0_n37_w118, 
            w119=> c0_n37_w119, 
            w120=> c0_n37_w120, 
            w121=> c0_n37_w121, 
            w122=> c0_n37_w122, 
            w123=> c0_n37_w123, 
            w124=> c0_n37_w124, 
            w125=> c0_n37_w125, 
            w126=> c0_n37_w126, 
            w127=> c0_n37_w127, 
            w128=> c0_n37_w128, 
            w129=> c0_n37_w129, 
            w130=> c0_n37_w130, 
            w131=> c0_n37_w131, 
            w132=> c0_n37_w132, 
            w133=> c0_n37_w133, 
            w134=> c0_n37_w134, 
            w135=> c0_n37_w135, 
            w136=> c0_n37_w136, 
            w137=> c0_n37_w137, 
            w138=> c0_n37_w138, 
            w139=> c0_n37_w139, 
            w140=> c0_n37_w140, 
            w141=> c0_n37_w141, 
            w142=> c0_n37_w142, 
            w143=> c0_n37_w143, 
            w144=> c0_n37_w144, 
            w145=> c0_n37_w145, 
            w146=> c0_n37_w146, 
            w147=> c0_n37_w147, 
            w148=> c0_n37_w148, 
            w149=> c0_n37_w149, 
            w150=> c0_n37_w150, 
            w151=> c0_n37_w151, 
            w152=> c0_n37_w152, 
            w153=> c0_n37_w153, 
            w154=> c0_n37_w154, 
            w155=> c0_n37_w155, 
            w156=> c0_n37_w156, 
            w157=> c0_n37_w157, 
            w158=> c0_n37_w158, 
            w159=> c0_n37_w159, 
            w160=> c0_n37_w160, 
            w161=> c0_n37_w161, 
            w162=> c0_n37_w162, 
            w163=> c0_n37_w163, 
            w164=> c0_n37_w164, 
            w165=> c0_n37_w165, 
            w166=> c0_n37_w166, 
            w167=> c0_n37_w167, 
            w168=> c0_n37_w168, 
            w169=> c0_n37_w169, 
            w170=> c0_n37_w170, 
            w171=> c0_n37_w171, 
            w172=> c0_n37_w172, 
            w173=> c0_n37_w173, 
            w174=> c0_n37_w174, 
            w175=> c0_n37_w175, 
            w176=> c0_n37_w176, 
            w177=> c0_n37_w177, 
            w178=> c0_n37_w178, 
            w179=> c0_n37_w179, 
            w180=> c0_n37_w180, 
            w181=> c0_n37_w181, 
            w182=> c0_n37_w182, 
            w183=> c0_n37_w183, 
            w184=> c0_n37_w184, 
            w185=> c0_n37_w185, 
            w186=> c0_n37_w186, 
            w187=> c0_n37_w187, 
            w188=> c0_n37_w188, 
            w189=> c0_n37_w189, 
            w190=> c0_n37_w190, 
            w191=> c0_n37_w191, 
            w192=> c0_n37_w192, 
            w193=> c0_n37_w193, 
            w194=> c0_n37_w194, 
            w195=> c0_n37_w195, 
            w196=> c0_n37_w196, 
            w197=> c0_n37_w197, 
            w198=> c0_n37_w198, 
            w199=> c0_n37_w199, 
            w200=> c0_n37_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n37_y
   );           
            
neuron_inst_38: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n38_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n38_w1, 
            w2=> c0_n38_w2, 
            w3=> c0_n38_w3, 
            w4=> c0_n38_w4, 
            w5=> c0_n38_w5, 
            w6=> c0_n38_w6, 
            w7=> c0_n38_w7, 
            w8=> c0_n38_w8, 
            w9=> c0_n38_w9, 
            w10=> c0_n38_w10, 
            w11=> c0_n38_w11, 
            w12=> c0_n38_w12, 
            w13=> c0_n38_w13, 
            w14=> c0_n38_w14, 
            w15=> c0_n38_w15, 
            w16=> c0_n38_w16, 
            w17=> c0_n38_w17, 
            w18=> c0_n38_w18, 
            w19=> c0_n38_w19, 
            w20=> c0_n38_w20, 
            w21=> c0_n38_w21, 
            w22=> c0_n38_w22, 
            w23=> c0_n38_w23, 
            w24=> c0_n38_w24, 
            w25=> c0_n38_w25, 
            w26=> c0_n38_w26, 
            w27=> c0_n38_w27, 
            w28=> c0_n38_w28, 
            w29=> c0_n38_w29, 
            w30=> c0_n38_w30, 
            w31=> c0_n38_w31, 
            w32=> c0_n38_w32, 
            w33=> c0_n38_w33, 
            w34=> c0_n38_w34, 
            w35=> c0_n38_w35, 
            w36=> c0_n38_w36, 
            w37=> c0_n38_w37, 
            w38=> c0_n38_w38, 
            w39=> c0_n38_w39, 
            w40=> c0_n38_w40, 
            w41=> c0_n38_w41, 
            w42=> c0_n38_w42, 
            w43=> c0_n38_w43, 
            w44=> c0_n38_w44, 
            w45=> c0_n38_w45, 
            w46=> c0_n38_w46, 
            w47=> c0_n38_w47, 
            w48=> c0_n38_w48, 
            w49=> c0_n38_w49, 
            w50=> c0_n38_w50, 
            w51=> c0_n38_w51, 
            w52=> c0_n38_w52, 
            w53=> c0_n38_w53, 
            w54=> c0_n38_w54, 
            w55=> c0_n38_w55, 
            w56=> c0_n38_w56, 
            w57=> c0_n38_w57, 
            w58=> c0_n38_w58, 
            w59=> c0_n38_w59, 
            w60=> c0_n38_w60, 
            w61=> c0_n38_w61, 
            w62=> c0_n38_w62, 
            w63=> c0_n38_w63, 
            w64=> c0_n38_w64, 
            w65=> c0_n38_w65, 
            w66=> c0_n38_w66, 
            w67=> c0_n38_w67, 
            w68=> c0_n38_w68, 
            w69=> c0_n38_w69, 
            w70=> c0_n38_w70, 
            w71=> c0_n38_w71, 
            w72=> c0_n38_w72, 
            w73=> c0_n38_w73, 
            w74=> c0_n38_w74, 
            w75=> c0_n38_w75, 
            w76=> c0_n38_w76, 
            w77=> c0_n38_w77, 
            w78=> c0_n38_w78, 
            w79=> c0_n38_w79, 
            w80=> c0_n38_w80, 
            w81=> c0_n38_w81, 
            w82=> c0_n38_w82, 
            w83=> c0_n38_w83, 
            w84=> c0_n38_w84, 
            w85=> c0_n38_w85, 
            w86=> c0_n38_w86, 
            w87=> c0_n38_w87, 
            w88=> c0_n38_w88, 
            w89=> c0_n38_w89, 
            w90=> c0_n38_w90, 
            w91=> c0_n38_w91, 
            w92=> c0_n38_w92, 
            w93=> c0_n38_w93, 
            w94=> c0_n38_w94, 
            w95=> c0_n38_w95, 
            w96=> c0_n38_w96, 
            w97=> c0_n38_w97, 
            w98=> c0_n38_w98, 
            w99=> c0_n38_w99, 
            w100=> c0_n38_w100, 
            w101=> c0_n38_w101, 
            w102=> c0_n38_w102, 
            w103=> c0_n38_w103, 
            w104=> c0_n38_w104, 
            w105=> c0_n38_w105, 
            w106=> c0_n38_w106, 
            w107=> c0_n38_w107, 
            w108=> c0_n38_w108, 
            w109=> c0_n38_w109, 
            w110=> c0_n38_w110, 
            w111=> c0_n38_w111, 
            w112=> c0_n38_w112, 
            w113=> c0_n38_w113, 
            w114=> c0_n38_w114, 
            w115=> c0_n38_w115, 
            w116=> c0_n38_w116, 
            w117=> c0_n38_w117, 
            w118=> c0_n38_w118, 
            w119=> c0_n38_w119, 
            w120=> c0_n38_w120, 
            w121=> c0_n38_w121, 
            w122=> c0_n38_w122, 
            w123=> c0_n38_w123, 
            w124=> c0_n38_w124, 
            w125=> c0_n38_w125, 
            w126=> c0_n38_w126, 
            w127=> c0_n38_w127, 
            w128=> c0_n38_w128, 
            w129=> c0_n38_w129, 
            w130=> c0_n38_w130, 
            w131=> c0_n38_w131, 
            w132=> c0_n38_w132, 
            w133=> c0_n38_w133, 
            w134=> c0_n38_w134, 
            w135=> c0_n38_w135, 
            w136=> c0_n38_w136, 
            w137=> c0_n38_w137, 
            w138=> c0_n38_w138, 
            w139=> c0_n38_w139, 
            w140=> c0_n38_w140, 
            w141=> c0_n38_w141, 
            w142=> c0_n38_w142, 
            w143=> c0_n38_w143, 
            w144=> c0_n38_w144, 
            w145=> c0_n38_w145, 
            w146=> c0_n38_w146, 
            w147=> c0_n38_w147, 
            w148=> c0_n38_w148, 
            w149=> c0_n38_w149, 
            w150=> c0_n38_w150, 
            w151=> c0_n38_w151, 
            w152=> c0_n38_w152, 
            w153=> c0_n38_w153, 
            w154=> c0_n38_w154, 
            w155=> c0_n38_w155, 
            w156=> c0_n38_w156, 
            w157=> c0_n38_w157, 
            w158=> c0_n38_w158, 
            w159=> c0_n38_w159, 
            w160=> c0_n38_w160, 
            w161=> c0_n38_w161, 
            w162=> c0_n38_w162, 
            w163=> c0_n38_w163, 
            w164=> c0_n38_w164, 
            w165=> c0_n38_w165, 
            w166=> c0_n38_w166, 
            w167=> c0_n38_w167, 
            w168=> c0_n38_w168, 
            w169=> c0_n38_w169, 
            w170=> c0_n38_w170, 
            w171=> c0_n38_w171, 
            w172=> c0_n38_w172, 
            w173=> c0_n38_w173, 
            w174=> c0_n38_w174, 
            w175=> c0_n38_w175, 
            w176=> c0_n38_w176, 
            w177=> c0_n38_w177, 
            w178=> c0_n38_w178, 
            w179=> c0_n38_w179, 
            w180=> c0_n38_w180, 
            w181=> c0_n38_w181, 
            w182=> c0_n38_w182, 
            w183=> c0_n38_w183, 
            w184=> c0_n38_w184, 
            w185=> c0_n38_w185, 
            w186=> c0_n38_w186, 
            w187=> c0_n38_w187, 
            w188=> c0_n38_w188, 
            w189=> c0_n38_w189, 
            w190=> c0_n38_w190, 
            w191=> c0_n38_w191, 
            w192=> c0_n38_w192, 
            w193=> c0_n38_w193, 
            w194=> c0_n38_w194, 
            w195=> c0_n38_w195, 
            w196=> c0_n38_w196, 
            w197=> c0_n38_w197, 
            w198=> c0_n38_w198, 
            w199=> c0_n38_w199, 
            w200=> c0_n38_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n38_y
   );           
            
neuron_inst_39: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n39_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n39_w1, 
            w2=> c0_n39_w2, 
            w3=> c0_n39_w3, 
            w4=> c0_n39_w4, 
            w5=> c0_n39_w5, 
            w6=> c0_n39_w6, 
            w7=> c0_n39_w7, 
            w8=> c0_n39_w8, 
            w9=> c0_n39_w9, 
            w10=> c0_n39_w10, 
            w11=> c0_n39_w11, 
            w12=> c0_n39_w12, 
            w13=> c0_n39_w13, 
            w14=> c0_n39_w14, 
            w15=> c0_n39_w15, 
            w16=> c0_n39_w16, 
            w17=> c0_n39_w17, 
            w18=> c0_n39_w18, 
            w19=> c0_n39_w19, 
            w20=> c0_n39_w20, 
            w21=> c0_n39_w21, 
            w22=> c0_n39_w22, 
            w23=> c0_n39_w23, 
            w24=> c0_n39_w24, 
            w25=> c0_n39_w25, 
            w26=> c0_n39_w26, 
            w27=> c0_n39_w27, 
            w28=> c0_n39_w28, 
            w29=> c0_n39_w29, 
            w30=> c0_n39_w30, 
            w31=> c0_n39_w31, 
            w32=> c0_n39_w32, 
            w33=> c0_n39_w33, 
            w34=> c0_n39_w34, 
            w35=> c0_n39_w35, 
            w36=> c0_n39_w36, 
            w37=> c0_n39_w37, 
            w38=> c0_n39_w38, 
            w39=> c0_n39_w39, 
            w40=> c0_n39_w40, 
            w41=> c0_n39_w41, 
            w42=> c0_n39_w42, 
            w43=> c0_n39_w43, 
            w44=> c0_n39_w44, 
            w45=> c0_n39_w45, 
            w46=> c0_n39_w46, 
            w47=> c0_n39_w47, 
            w48=> c0_n39_w48, 
            w49=> c0_n39_w49, 
            w50=> c0_n39_w50, 
            w51=> c0_n39_w51, 
            w52=> c0_n39_w52, 
            w53=> c0_n39_w53, 
            w54=> c0_n39_w54, 
            w55=> c0_n39_w55, 
            w56=> c0_n39_w56, 
            w57=> c0_n39_w57, 
            w58=> c0_n39_w58, 
            w59=> c0_n39_w59, 
            w60=> c0_n39_w60, 
            w61=> c0_n39_w61, 
            w62=> c0_n39_w62, 
            w63=> c0_n39_w63, 
            w64=> c0_n39_w64, 
            w65=> c0_n39_w65, 
            w66=> c0_n39_w66, 
            w67=> c0_n39_w67, 
            w68=> c0_n39_w68, 
            w69=> c0_n39_w69, 
            w70=> c0_n39_w70, 
            w71=> c0_n39_w71, 
            w72=> c0_n39_w72, 
            w73=> c0_n39_w73, 
            w74=> c0_n39_w74, 
            w75=> c0_n39_w75, 
            w76=> c0_n39_w76, 
            w77=> c0_n39_w77, 
            w78=> c0_n39_w78, 
            w79=> c0_n39_w79, 
            w80=> c0_n39_w80, 
            w81=> c0_n39_w81, 
            w82=> c0_n39_w82, 
            w83=> c0_n39_w83, 
            w84=> c0_n39_w84, 
            w85=> c0_n39_w85, 
            w86=> c0_n39_w86, 
            w87=> c0_n39_w87, 
            w88=> c0_n39_w88, 
            w89=> c0_n39_w89, 
            w90=> c0_n39_w90, 
            w91=> c0_n39_w91, 
            w92=> c0_n39_w92, 
            w93=> c0_n39_w93, 
            w94=> c0_n39_w94, 
            w95=> c0_n39_w95, 
            w96=> c0_n39_w96, 
            w97=> c0_n39_w97, 
            w98=> c0_n39_w98, 
            w99=> c0_n39_w99, 
            w100=> c0_n39_w100, 
            w101=> c0_n39_w101, 
            w102=> c0_n39_w102, 
            w103=> c0_n39_w103, 
            w104=> c0_n39_w104, 
            w105=> c0_n39_w105, 
            w106=> c0_n39_w106, 
            w107=> c0_n39_w107, 
            w108=> c0_n39_w108, 
            w109=> c0_n39_w109, 
            w110=> c0_n39_w110, 
            w111=> c0_n39_w111, 
            w112=> c0_n39_w112, 
            w113=> c0_n39_w113, 
            w114=> c0_n39_w114, 
            w115=> c0_n39_w115, 
            w116=> c0_n39_w116, 
            w117=> c0_n39_w117, 
            w118=> c0_n39_w118, 
            w119=> c0_n39_w119, 
            w120=> c0_n39_w120, 
            w121=> c0_n39_w121, 
            w122=> c0_n39_w122, 
            w123=> c0_n39_w123, 
            w124=> c0_n39_w124, 
            w125=> c0_n39_w125, 
            w126=> c0_n39_w126, 
            w127=> c0_n39_w127, 
            w128=> c0_n39_w128, 
            w129=> c0_n39_w129, 
            w130=> c0_n39_w130, 
            w131=> c0_n39_w131, 
            w132=> c0_n39_w132, 
            w133=> c0_n39_w133, 
            w134=> c0_n39_w134, 
            w135=> c0_n39_w135, 
            w136=> c0_n39_w136, 
            w137=> c0_n39_w137, 
            w138=> c0_n39_w138, 
            w139=> c0_n39_w139, 
            w140=> c0_n39_w140, 
            w141=> c0_n39_w141, 
            w142=> c0_n39_w142, 
            w143=> c0_n39_w143, 
            w144=> c0_n39_w144, 
            w145=> c0_n39_w145, 
            w146=> c0_n39_w146, 
            w147=> c0_n39_w147, 
            w148=> c0_n39_w148, 
            w149=> c0_n39_w149, 
            w150=> c0_n39_w150, 
            w151=> c0_n39_w151, 
            w152=> c0_n39_w152, 
            w153=> c0_n39_w153, 
            w154=> c0_n39_w154, 
            w155=> c0_n39_w155, 
            w156=> c0_n39_w156, 
            w157=> c0_n39_w157, 
            w158=> c0_n39_w158, 
            w159=> c0_n39_w159, 
            w160=> c0_n39_w160, 
            w161=> c0_n39_w161, 
            w162=> c0_n39_w162, 
            w163=> c0_n39_w163, 
            w164=> c0_n39_w164, 
            w165=> c0_n39_w165, 
            w166=> c0_n39_w166, 
            w167=> c0_n39_w167, 
            w168=> c0_n39_w168, 
            w169=> c0_n39_w169, 
            w170=> c0_n39_w170, 
            w171=> c0_n39_w171, 
            w172=> c0_n39_w172, 
            w173=> c0_n39_w173, 
            w174=> c0_n39_w174, 
            w175=> c0_n39_w175, 
            w176=> c0_n39_w176, 
            w177=> c0_n39_w177, 
            w178=> c0_n39_w178, 
            w179=> c0_n39_w179, 
            w180=> c0_n39_w180, 
            w181=> c0_n39_w181, 
            w182=> c0_n39_w182, 
            w183=> c0_n39_w183, 
            w184=> c0_n39_w184, 
            w185=> c0_n39_w185, 
            w186=> c0_n39_w186, 
            w187=> c0_n39_w187, 
            w188=> c0_n39_w188, 
            w189=> c0_n39_w189, 
            w190=> c0_n39_w190, 
            w191=> c0_n39_w191, 
            w192=> c0_n39_w192, 
            w193=> c0_n39_w193, 
            w194=> c0_n39_w194, 
            w195=> c0_n39_w195, 
            w196=> c0_n39_w196, 
            w197=> c0_n39_w197, 
            w198=> c0_n39_w198, 
            w199=> c0_n39_w199, 
            w200=> c0_n39_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n39_y
   );           
            
neuron_inst_40: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n40_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n40_w1, 
            w2=> c0_n40_w2, 
            w3=> c0_n40_w3, 
            w4=> c0_n40_w4, 
            w5=> c0_n40_w5, 
            w6=> c0_n40_w6, 
            w7=> c0_n40_w7, 
            w8=> c0_n40_w8, 
            w9=> c0_n40_w9, 
            w10=> c0_n40_w10, 
            w11=> c0_n40_w11, 
            w12=> c0_n40_w12, 
            w13=> c0_n40_w13, 
            w14=> c0_n40_w14, 
            w15=> c0_n40_w15, 
            w16=> c0_n40_w16, 
            w17=> c0_n40_w17, 
            w18=> c0_n40_w18, 
            w19=> c0_n40_w19, 
            w20=> c0_n40_w20, 
            w21=> c0_n40_w21, 
            w22=> c0_n40_w22, 
            w23=> c0_n40_w23, 
            w24=> c0_n40_w24, 
            w25=> c0_n40_w25, 
            w26=> c0_n40_w26, 
            w27=> c0_n40_w27, 
            w28=> c0_n40_w28, 
            w29=> c0_n40_w29, 
            w30=> c0_n40_w30, 
            w31=> c0_n40_w31, 
            w32=> c0_n40_w32, 
            w33=> c0_n40_w33, 
            w34=> c0_n40_w34, 
            w35=> c0_n40_w35, 
            w36=> c0_n40_w36, 
            w37=> c0_n40_w37, 
            w38=> c0_n40_w38, 
            w39=> c0_n40_w39, 
            w40=> c0_n40_w40, 
            w41=> c0_n40_w41, 
            w42=> c0_n40_w42, 
            w43=> c0_n40_w43, 
            w44=> c0_n40_w44, 
            w45=> c0_n40_w45, 
            w46=> c0_n40_w46, 
            w47=> c0_n40_w47, 
            w48=> c0_n40_w48, 
            w49=> c0_n40_w49, 
            w50=> c0_n40_w50, 
            w51=> c0_n40_w51, 
            w52=> c0_n40_w52, 
            w53=> c0_n40_w53, 
            w54=> c0_n40_w54, 
            w55=> c0_n40_w55, 
            w56=> c0_n40_w56, 
            w57=> c0_n40_w57, 
            w58=> c0_n40_w58, 
            w59=> c0_n40_w59, 
            w60=> c0_n40_w60, 
            w61=> c0_n40_w61, 
            w62=> c0_n40_w62, 
            w63=> c0_n40_w63, 
            w64=> c0_n40_w64, 
            w65=> c0_n40_w65, 
            w66=> c0_n40_w66, 
            w67=> c0_n40_w67, 
            w68=> c0_n40_w68, 
            w69=> c0_n40_w69, 
            w70=> c0_n40_w70, 
            w71=> c0_n40_w71, 
            w72=> c0_n40_w72, 
            w73=> c0_n40_w73, 
            w74=> c0_n40_w74, 
            w75=> c0_n40_w75, 
            w76=> c0_n40_w76, 
            w77=> c0_n40_w77, 
            w78=> c0_n40_w78, 
            w79=> c0_n40_w79, 
            w80=> c0_n40_w80, 
            w81=> c0_n40_w81, 
            w82=> c0_n40_w82, 
            w83=> c0_n40_w83, 
            w84=> c0_n40_w84, 
            w85=> c0_n40_w85, 
            w86=> c0_n40_w86, 
            w87=> c0_n40_w87, 
            w88=> c0_n40_w88, 
            w89=> c0_n40_w89, 
            w90=> c0_n40_w90, 
            w91=> c0_n40_w91, 
            w92=> c0_n40_w92, 
            w93=> c0_n40_w93, 
            w94=> c0_n40_w94, 
            w95=> c0_n40_w95, 
            w96=> c0_n40_w96, 
            w97=> c0_n40_w97, 
            w98=> c0_n40_w98, 
            w99=> c0_n40_w99, 
            w100=> c0_n40_w100, 
            w101=> c0_n40_w101, 
            w102=> c0_n40_w102, 
            w103=> c0_n40_w103, 
            w104=> c0_n40_w104, 
            w105=> c0_n40_w105, 
            w106=> c0_n40_w106, 
            w107=> c0_n40_w107, 
            w108=> c0_n40_w108, 
            w109=> c0_n40_w109, 
            w110=> c0_n40_w110, 
            w111=> c0_n40_w111, 
            w112=> c0_n40_w112, 
            w113=> c0_n40_w113, 
            w114=> c0_n40_w114, 
            w115=> c0_n40_w115, 
            w116=> c0_n40_w116, 
            w117=> c0_n40_w117, 
            w118=> c0_n40_w118, 
            w119=> c0_n40_w119, 
            w120=> c0_n40_w120, 
            w121=> c0_n40_w121, 
            w122=> c0_n40_w122, 
            w123=> c0_n40_w123, 
            w124=> c0_n40_w124, 
            w125=> c0_n40_w125, 
            w126=> c0_n40_w126, 
            w127=> c0_n40_w127, 
            w128=> c0_n40_w128, 
            w129=> c0_n40_w129, 
            w130=> c0_n40_w130, 
            w131=> c0_n40_w131, 
            w132=> c0_n40_w132, 
            w133=> c0_n40_w133, 
            w134=> c0_n40_w134, 
            w135=> c0_n40_w135, 
            w136=> c0_n40_w136, 
            w137=> c0_n40_w137, 
            w138=> c0_n40_w138, 
            w139=> c0_n40_w139, 
            w140=> c0_n40_w140, 
            w141=> c0_n40_w141, 
            w142=> c0_n40_w142, 
            w143=> c0_n40_w143, 
            w144=> c0_n40_w144, 
            w145=> c0_n40_w145, 
            w146=> c0_n40_w146, 
            w147=> c0_n40_w147, 
            w148=> c0_n40_w148, 
            w149=> c0_n40_w149, 
            w150=> c0_n40_w150, 
            w151=> c0_n40_w151, 
            w152=> c0_n40_w152, 
            w153=> c0_n40_w153, 
            w154=> c0_n40_w154, 
            w155=> c0_n40_w155, 
            w156=> c0_n40_w156, 
            w157=> c0_n40_w157, 
            w158=> c0_n40_w158, 
            w159=> c0_n40_w159, 
            w160=> c0_n40_w160, 
            w161=> c0_n40_w161, 
            w162=> c0_n40_w162, 
            w163=> c0_n40_w163, 
            w164=> c0_n40_w164, 
            w165=> c0_n40_w165, 
            w166=> c0_n40_w166, 
            w167=> c0_n40_w167, 
            w168=> c0_n40_w168, 
            w169=> c0_n40_w169, 
            w170=> c0_n40_w170, 
            w171=> c0_n40_w171, 
            w172=> c0_n40_w172, 
            w173=> c0_n40_w173, 
            w174=> c0_n40_w174, 
            w175=> c0_n40_w175, 
            w176=> c0_n40_w176, 
            w177=> c0_n40_w177, 
            w178=> c0_n40_w178, 
            w179=> c0_n40_w179, 
            w180=> c0_n40_w180, 
            w181=> c0_n40_w181, 
            w182=> c0_n40_w182, 
            w183=> c0_n40_w183, 
            w184=> c0_n40_w184, 
            w185=> c0_n40_w185, 
            w186=> c0_n40_w186, 
            w187=> c0_n40_w187, 
            w188=> c0_n40_w188, 
            w189=> c0_n40_w189, 
            w190=> c0_n40_w190, 
            w191=> c0_n40_w191, 
            w192=> c0_n40_w192, 
            w193=> c0_n40_w193, 
            w194=> c0_n40_w194, 
            w195=> c0_n40_w195, 
            w196=> c0_n40_w196, 
            w197=> c0_n40_w197, 
            w198=> c0_n40_w198, 
            w199=> c0_n40_w199, 
            w200=> c0_n40_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n40_y
   );           
            
neuron_inst_41: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n41_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n41_w1, 
            w2=> c0_n41_w2, 
            w3=> c0_n41_w3, 
            w4=> c0_n41_w4, 
            w5=> c0_n41_w5, 
            w6=> c0_n41_w6, 
            w7=> c0_n41_w7, 
            w8=> c0_n41_w8, 
            w9=> c0_n41_w9, 
            w10=> c0_n41_w10, 
            w11=> c0_n41_w11, 
            w12=> c0_n41_w12, 
            w13=> c0_n41_w13, 
            w14=> c0_n41_w14, 
            w15=> c0_n41_w15, 
            w16=> c0_n41_w16, 
            w17=> c0_n41_w17, 
            w18=> c0_n41_w18, 
            w19=> c0_n41_w19, 
            w20=> c0_n41_w20, 
            w21=> c0_n41_w21, 
            w22=> c0_n41_w22, 
            w23=> c0_n41_w23, 
            w24=> c0_n41_w24, 
            w25=> c0_n41_w25, 
            w26=> c0_n41_w26, 
            w27=> c0_n41_w27, 
            w28=> c0_n41_w28, 
            w29=> c0_n41_w29, 
            w30=> c0_n41_w30, 
            w31=> c0_n41_w31, 
            w32=> c0_n41_w32, 
            w33=> c0_n41_w33, 
            w34=> c0_n41_w34, 
            w35=> c0_n41_w35, 
            w36=> c0_n41_w36, 
            w37=> c0_n41_w37, 
            w38=> c0_n41_w38, 
            w39=> c0_n41_w39, 
            w40=> c0_n41_w40, 
            w41=> c0_n41_w41, 
            w42=> c0_n41_w42, 
            w43=> c0_n41_w43, 
            w44=> c0_n41_w44, 
            w45=> c0_n41_w45, 
            w46=> c0_n41_w46, 
            w47=> c0_n41_w47, 
            w48=> c0_n41_w48, 
            w49=> c0_n41_w49, 
            w50=> c0_n41_w50, 
            w51=> c0_n41_w51, 
            w52=> c0_n41_w52, 
            w53=> c0_n41_w53, 
            w54=> c0_n41_w54, 
            w55=> c0_n41_w55, 
            w56=> c0_n41_w56, 
            w57=> c0_n41_w57, 
            w58=> c0_n41_w58, 
            w59=> c0_n41_w59, 
            w60=> c0_n41_w60, 
            w61=> c0_n41_w61, 
            w62=> c0_n41_w62, 
            w63=> c0_n41_w63, 
            w64=> c0_n41_w64, 
            w65=> c0_n41_w65, 
            w66=> c0_n41_w66, 
            w67=> c0_n41_w67, 
            w68=> c0_n41_w68, 
            w69=> c0_n41_w69, 
            w70=> c0_n41_w70, 
            w71=> c0_n41_w71, 
            w72=> c0_n41_w72, 
            w73=> c0_n41_w73, 
            w74=> c0_n41_w74, 
            w75=> c0_n41_w75, 
            w76=> c0_n41_w76, 
            w77=> c0_n41_w77, 
            w78=> c0_n41_w78, 
            w79=> c0_n41_w79, 
            w80=> c0_n41_w80, 
            w81=> c0_n41_w81, 
            w82=> c0_n41_w82, 
            w83=> c0_n41_w83, 
            w84=> c0_n41_w84, 
            w85=> c0_n41_w85, 
            w86=> c0_n41_w86, 
            w87=> c0_n41_w87, 
            w88=> c0_n41_w88, 
            w89=> c0_n41_w89, 
            w90=> c0_n41_w90, 
            w91=> c0_n41_w91, 
            w92=> c0_n41_w92, 
            w93=> c0_n41_w93, 
            w94=> c0_n41_w94, 
            w95=> c0_n41_w95, 
            w96=> c0_n41_w96, 
            w97=> c0_n41_w97, 
            w98=> c0_n41_w98, 
            w99=> c0_n41_w99, 
            w100=> c0_n41_w100, 
            w101=> c0_n41_w101, 
            w102=> c0_n41_w102, 
            w103=> c0_n41_w103, 
            w104=> c0_n41_w104, 
            w105=> c0_n41_w105, 
            w106=> c0_n41_w106, 
            w107=> c0_n41_w107, 
            w108=> c0_n41_w108, 
            w109=> c0_n41_w109, 
            w110=> c0_n41_w110, 
            w111=> c0_n41_w111, 
            w112=> c0_n41_w112, 
            w113=> c0_n41_w113, 
            w114=> c0_n41_w114, 
            w115=> c0_n41_w115, 
            w116=> c0_n41_w116, 
            w117=> c0_n41_w117, 
            w118=> c0_n41_w118, 
            w119=> c0_n41_w119, 
            w120=> c0_n41_w120, 
            w121=> c0_n41_w121, 
            w122=> c0_n41_w122, 
            w123=> c0_n41_w123, 
            w124=> c0_n41_w124, 
            w125=> c0_n41_w125, 
            w126=> c0_n41_w126, 
            w127=> c0_n41_w127, 
            w128=> c0_n41_w128, 
            w129=> c0_n41_w129, 
            w130=> c0_n41_w130, 
            w131=> c0_n41_w131, 
            w132=> c0_n41_w132, 
            w133=> c0_n41_w133, 
            w134=> c0_n41_w134, 
            w135=> c0_n41_w135, 
            w136=> c0_n41_w136, 
            w137=> c0_n41_w137, 
            w138=> c0_n41_w138, 
            w139=> c0_n41_w139, 
            w140=> c0_n41_w140, 
            w141=> c0_n41_w141, 
            w142=> c0_n41_w142, 
            w143=> c0_n41_w143, 
            w144=> c0_n41_w144, 
            w145=> c0_n41_w145, 
            w146=> c0_n41_w146, 
            w147=> c0_n41_w147, 
            w148=> c0_n41_w148, 
            w149=> c0_n41_w149, 
            w150=> c0_n41_w150, 
            w151=> c0_n41_w151, 
            w152=> c0_n41_w152, 
            w153=> c0_n41_w153, 
            w154=> c0_n41_w154, 
            w155=> c0_n41_w155, 
            w156=> c0_n41_w156, 
            w157=> c0_n41_w157, 
            w158=> c0_n41_w158, 
            w159=> c0_n41_w159, 
            w160=> c0_n41_w160, 
            w161=> c0_n41_w161, 
            w162=> c0_n41_w162, 
            w163=> c0_n41_w163, 
            w164=> c0_n41_w164, 
            w165=> c0_n41_w165, 
            w166=> c0_n41_w166, 
            w167=> c0_n41_w167, 
            w168=> c0_n41_w168, 
            w169=> c0_n41_w169, 
            w170=> c0_n41_w170, 
            w171=> c0_n41_w171, 
            w172=> c0_n41_w172, 
            w173=> c0_n41_w173, 
            w174=> c0_n41_w174, 
            w175=> c0_n41_w175, 
            w176=> c0_n41_w176, 
            w177=> c0_n41_w177, 
            w178=> c0_n41_w178, 
            w179=> c0_n41_w179, 
            w180=> c0_n41_w180, 
            w181=> c0_n41_w181, 
            w182=> c0_n41_w182, 
            w183=> c0_n41_w183, 
            w184=> c0_n41_w184, 
            w185=> c0_n41_w185, 
            w186=> c0_n41_w186, 
            w187=> c0_n41_w187, 
            w188=> c0_n41_w188, 
            w189=> c0_n41_w189, 
            w190=> c0_n41_w190, 
            w191=> c0_n41_w191, 
            w192=> c0_n41_w192, 
            w193=> c0_n41_w193, 
            w194=> c0_n41_w194, 
            w195=> c0_n41_w195, 
            w196=> c0_n41_w196, 
            w197=> c0_n41_w197, 
            w198=> c0_n41_w198, 
            w199=> c0_n41_w199, 
            w200=> c0_n41_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n41_y
   );           
            
neuron_inst_42: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n42_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n42_w1, 
            w2=> c0_n42_w2, 
            w3=> c0_n42_w3, 
            w4=> c0_n42_w4, 
            w5=> c0_n42_w5, 
            w6=> c0_n42_w6, 
            w7=> c0_n42_w7, 
            w8=> c0_n42_w8, 
            w9=> c0_n42_w9, 
            w10=> c0_n42_w10, 
            w11=> c0_n42_w11, 
            w12=> c0_n42_w12, 
            w13=> c0_n42_w13, 
            w14=> c0_n42_w14, 
            w15=> c0_n42_w15, 
            w16=> c0_n42_w16, 
            w17=> c0_n42_w17, 
            w18=> c0_n42_w18, 
            w19=> c0_n42_w19, 
            w20=> c0_n42_w20, 
            w21=> c0_n42_w21, 
            w22=> c0_n42_w22, 
            w23=> c0_n42_w23, 
            w24=> c0_n42_w24, 
            w25=> c0_n42_w25, 
            w26=> c0_n42_w26, 
            w27=> c0_n42_w27, 
            w28=> c0_n42_w28, 
            w29=> c0_n42_w29, 
            w30=> c0_n42_w30, 
            w31=> c0_n42_w31, 
            w32=> c0_n42_w32, 
            w33=> c0_n42_w33, 
            w34=> c0_n42_w34, 
            w35=> c0_n42_w35, 
            w36=> c0_n42_w36, 
            w37=> c0_n42_w37, 
            w38=> c0_n42_w38, 
            w39=> c0_n42_w39, 
            w40=> c0_n42_w40, 
            w41=> c0_n42_w41, 
            w42=> c0_n42_w42, 
            w43=> c0_n42_w43, 
            w44=> c0_n42_w44, 
            w45=> c0_n42_w45, 
            w46=> c0_n42_w46, 
            w47=> c0_n42_w47, 
            w48=> c0_n42_w48, 
            w49=> c0_n42_w49, 
            w50=> c0_n42_w50, 
            w51=> c0_n42_w51, 
            w52=> c0_n42_w52, 
            w53=> c0_n42_w53, 
            w54=> c0_n42_w54, 
            w55=> c0_n42_w55, 
            w56=> c0_n42_w56, 
            w57=> c0_n42_w57, 
            w58=> c0_n42_w58, 
            w59=> c0_n42_w59, 
            w60=> c0_n42_w60, 
            w61=> c0_n42_w61, 
            w62=> c0_n42_w62, 
            w63=> c0_n42_w63, 
            w64=> c0_n42_w64, 
            w65=> c0_n42_w65, 
            w66=> c0_n42_w66, 
            w67=> c0_n42_w67, 
            w68=> c0_n42_w68, 
            w69=> c0_n42_w69, 
            w70=> c0_n42_w70, 
            w71=> c0_n42_w71, 
            w72=> c0_n42_w72, 
            w73=> c0_n42_w73, 
            w74=> c0_n42_w74, 
            w75=> c0_n42_w75, 
            w76=> c0_n42_w76, 
            w77=> c0_n42_w77, 
            w78=> c0_n42_w78, 
            w79=> c0_n42_w79, 
            w80=> c0_n42_w80, 
            w81=> c0_n42_w81, 
            w82=> c0_n42_w82, 
            w83=> c0_n42_w83, 
            w84=> c0_n42_w84, 
            w85=> c0_n42_w85, 
            w86=> c0_n42_w86, 
            w87=> c0_n42_w87, 
            w88=> c0_n42_w88, 
            w89=> c0_n42_w89, 
            w90=> c0_n42_w90, 
            w91=> c0_n42_w91, 
            w92=> c0_n42_w92, 
            w93=> c0_n42_w93, 
            w94=> c0_n42_w94, 
            w95=> c0_n42_w95, 
            w96=> c0_n42_w96, 
            w97=> c0_n42_w97, 
            w98=> c0_n42_w98, 
            w99=> c0_n42_w99, 
            w100=> c0_n42_w100, 
            w101=> c0_n42_w101, 
            w102=> c0_n42_w102, 
            w103=> c0_n42_w103, 
            w104=> c0_n42_w104, 
            w105=> c0_n42_w105, 
            w106=> c0_n42_w106, 
            w107=> c0_n42_w107, 
            w108=> c0_n42_w108, 
            w109=> c0_n42_w109, 
            w110=> c0_n42_w110, 
            w111=> c0_n42_w111, 
            w112=> c0_n42_w112, 
            w113=> c0_n42_w113, 
            w114=> c0_n42_w114, 
            w115=> c0_n42_w115, 
            w116=> c0_n42_w116, 
            w117=> c0_n42_w117, 
            w118=> c0_n42_w118, 
            w119=> c0_n42_w119, 
            w120=> c0_n42_w120, 
            w121=> c0_n42_w121, 
            w122=> c0_n42_w122, 
            w123=> c0_n42_w123, 
            w124=> c0_n42_w124, 
            w125=> c0_n42_w125, 
            w126=> c0_n42_w126, 
            w127=> c0_n42_w127, 
            w128=> c0_n42_w128, 
            w129=> c0_n42_w129, 
            w130=> c0_n42_w130, 
            w131=> c0_n42_w131, 
            w132=> c0_n42_w132, 
            w133=> c0_n42_w133, 
            w134=> c0_n42_w134, 
            w135=> c0_n42_w135, 
            w136=> c0_n42_w136, 
            w137=> c0_n42_w137, 
            w138=> c0_n42_w138, 
            w139=> c0_n42_w139, 
            w140=> c0_n42_w140, 
            w141=> c0_n42_w141, 
            w142=> c0_n42_w142, 
            w143=> c0_n42_w143, 
            w144=> c0_n42_w144, 
            w145=> c0_n42_w145, 
            w146=> c0_n42_w146, 
            w147=> c0_n42_w147, 
            w148=> c0_n42_w148, 
            w149=> c0_n42_w149, 
            w150=> c0_n42_w150, 
            w151=> c0_n42_w151, 
            w152=> c0_n42_w152, 
            w153=> c0_n42_w153, 
            w154=> c0_n42_w154, 
            w155=> c0_n42_w155, 
            w156=> c0_n42_w156, 
            w157=> c0_n42_w157, 
            w158=> c0_n42_w158, 
            w159=> c0_n42_w159, 
            w160=> c0_n42_w160, 
            w161=> c0_n42_w161, 
            w162=> c0_n42_w162, 
            w163=> c0_n42_w163, 
            w164=> c0_n42_w164, 
            w165=> c0_n42_w165, 
            w166=> c0_n42_w166, 
            w167=> c0_n42_w167, 
            w168=> c0_n42_w168, 
            w169=> c0_n42_w169, 
            w170=> c0_n42_w170, 
            w171=> c0_n42_w171, 
            w172=> c0_n42_w172, 
            w173=> c0_n42_w173, 
            w174=> c0_n42_w174, 
            w175=> c0_n42_w175, 
            w176=> c0_n42_w176, 
            w177=> c0_n42_w177, 
            w178=> c0_n42_w178, 
            w179=> c0_n42_w179, 
            w180=> c0_n42_w180, 
            w181=> c0_n42_w181, 
            w182=> c0_n42_w182, 
            w183=> c0_n42_w183, 
            w184=> c0_n42_w184, 
            w185=> c0_n42_w185, 
            w186=> c0_n42_w186, 
            w187=> c0_n42_w187, 
            w188=> c0_n42_w188, 
            w189=> c0_n42_w189, 
            w190=> c0_n42_w190, 
            w191=> c0_n42_w191, 
            w192=> c0_n42_w192, 
            w193=> c0_n42_w193, 
            w194=> c0_n42_w194, 
            w195=> c0_n42_w195, 
            w196=> c0_n42_w196, 
            w197=> c0_n42_w197, 
            w198=> c0_n42_w198, 
            w199=> c0_n42_w199, 
            w200=> c0_n42_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n42_y
   );           
            
neuron_inst_43: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n43_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n43_w1, 
            w2=> c0_n43_w2, 
            w3=> c0_n43_w3, 
            w4=> c0_n43_w4, 
            w5=> c0_n43_w5, 
            w6=> c0_n43_w6, 
            w7=> c0_n43_w7, 
            w8=> c0_n43_w8, 
            w9=> c0_n43_w9, 
            w10=> c0_n43_w10, 
            w11=> c0_n43_w11, 
            w12=> c0_n43_w12, 
            w13=> c0_n43_w13, 
            w14=> c0_n43_w14, 
            w15=> c0_n43_w15, 
            w16=> c0_n43_w16, 
            w17=> c0_n43_w17, 
            w18=> c0_n43_w18, 
            w19=> c0_n43_w19, 
            w20=> c0_n43_w20, 
            w21=> c0_n43_w21, 
            w22=> c0_n43_w22, 
            w23=> c0_n43_w23, 
            w24=> c0_n43_w24, 
            w25=> c0_n43_w25, 
            w26=> c0_n43_w26, 
            w27=> c0_n43_w27, 
            w28=> c0_n43_w28, 
            w29=> c0_n43_w29, 
            w30=> c0_n43_w30, 
            w31=> c0_n43_w31, 
            w32=> c0_n43_w32, 
            w33=> c0_n43_w33, 
            w34=> c0_n43_w34, 
            w35=> c0_n43_w35, 
            w36=> c0_n43_w36, 
            w37=> c0_n43_w37, 
            w38=> c0_n43_w38, 
            w39=> c0_n43_w39, 
            w40=> c0_n43_w40, 
            w41=> c0_n43_w41, 
            w42=> c0_n43_w42, 
            w43=> c0_n43_w43, 
            w44=> c0_n43_w44, 
            w45=> c0_n43_w45, 
            w46=> c0_n43_w46, 
            w47=> c0_n43_w47, 
            w48=> c0_n43_w48, 
            w49=> c0_n43_w49, 
            w50=> c0_n43_w50, 
            w51=> c0_n43_w51, 
            w52=> c0_n43_w52, 
            w53=> c0_n43_w53, 
            w54=> c0_n43_w54, 
            w55=> c0_n43_w55, 
            w56=> c0_n43_w56, 
            w57=> c0_n43_w57, 
            w58=> c0_n43_w58, 
            w59=> c0_n43_w59, 
            w60=> c0_n43_w60, 
            w61=> c0_n43_w61, 
            w62=> c0_n43_w62, 
            w63=> c0_n43_w63, 
            w64=> c0_n43_w64, 
            w65=> c0_n43_w65, 
            w66=> c0_n43_w66, 
            w67=> c0_n43_w67, 
            w68=> c0_n43_w68, 
            w69=> c0_n43_w69, 
            w70=> c0_n43_w70, 
            w71=> c0_n43_w71, 
            w72=> c0_n43_w72, 
            w73=> c0_n43_w73, 
            w74=> c0_n43_w74, 
            w75=> c0_n43_w75, 
            w76=> c0_n43_w76, 
            w77=> c0_n43_w77, 
            w78=> c0_n43_w78, 
            w79=> c0_n43_w79, 
            w80=> c0_n43_w80, 
            w81=> c0_n43_w81, 
            w82=> c0_n43_w82, 
            w83=> c0_n43_w83, 
            w84=> c0_n43_w84, 
            w85=> c0_n43_w85, 
            w86=> c0_n43_w86, 
            w87=> c0_n43_w87, 
            w88=> c0_n43_w88, 
            w89=> c0_n43_w89, 
            w90=> c0_n43_w90, 
            w91=> c0_n43_w91, 
            w92=> c0_n43_w92, 
            w93=> c0_n43_w93, 
            w94=> c0_n43_w94, 
            w95=> c0_n43_w95, 
            w96=> c0_n43_w96, 
            w97=> c0_n43_w97, 
            w98=> c0_n43_w98, 
            w99=> c0_n43_w99, 
            w100=> c0_n43_w100, 
            w101=> c0_n43_w101, 
            w102=> c0_n43_w102, 
            w103=> c0_n43_w103, 
            w104=> c0_n43_w104, 
            w105=> c0_n43_w105, 
            w106=> c0_n43_w106, 
            w107=> c0_n43_w107, 
            w108=> c0_n43_w108, 
            w109=> c0_n43_w109, 
            w110=> c0_n43_w110, 
            w111=> c0_n43_w111, 
            w112=> c0_n43_w112, 
            w113=> c0_n43_w113, 
            w114=> c0_n43_w114, 
            w115=> c0_n43_w115, 
            w116=> c0_n43_w116, 
            w117=> c0_n43_w117, 
            w118=> c0_n43_w118, 
            w119=> c0_n43_w119, 
            w120=> c0_n43_w120, 
            w121=> c0_n43_w121, 
            w122=> c0_n43_w122, 
            w123=> c0_n43_w123, 
            w124=> c0_n43_w124, 
            w125=> c0_n43_w125, 
            w126=> c0_n43_w126, 
            w127=> c0_n43_w127, 
            w128=> c0_n43_w128, 
            w129=> c0_n43_w129, 
            w130=> c0_n43_w130, 
            w131=> c0_n43_w131, 
            w132=> c0_n43_w132, 
            w133=> c0_n43_w133, 
            w134=> c0_n43_w134, 
            w135=> c0_n43_w135, 
            w136=> c0_n43_w136, 
            w137=> c0_n43_w137, 
            w138=> c0_n43_w138, 
            w139=> c0_n43_w139, 
            w140=> c0_n43_w140, 
            w141=> c0_n43_w141, 
            w142=> c0_n43_w142, 
            w143=> c0_n43_w143, 
            w144=> c0_n43_w144, 
            w145=> c0_n43_w145, 
            w146=> c0_n43_w146, 
            w147=> c0_n43_w147, 
            w148=> c0_n43_w148, 
            w149=> c0_n43_w149, 
            w150=> c0_n43_w150, 
            w151=> c0_n43_w151, 
            w152=> c0_n43_w152, 
            w153=> c0_n43_w153, 
            w154=> c0_n43_w154, 
            w155=> c0_n43_w155, 
            w156=> c0_n43_w156, 
            w157=> c0_n43_w157, 
            w158=> c0_n43_w158, 
            w159=> c0_n43_w159, 
            w160=> c0_n43_w160, 
            w161=> c0_n43_w161, 
            w162=> c0_n43_w162, 
            w163=> c0_n43_w163, 
            w164=> c0_n43_w164, 
            w165=> c0_n43_w165, 
            w166=> c0_n43_w166, 
            w167=> c0_n43_w167, 
            w168=> c0_n43_w168, 
            w169=> c0_n43_w169, 
            w170=> c0_n43_w170, 
            w171=> c0_n43_w171, 
            w172=> c0_n43_w172, 
            w173=> c0_n43_w173, 
            w174=> c0_n43_w174, 
            w175=> c0_n43_w175, 
            w176=> c0_n43_w176, 
            w177=> c0_n43_w177, 
            w178=> c0_n43_w178, 
            w179=> c0_n43_w179, 
            w180=> c0_n43_w180, 
            w181=> c0_n43_w181, 
            w182=> c0_n43_w182, 
            w183=> c0_n43_w183, 
            w184=> c0_n43_w184, 
            w185=> c0_n43_w185, 
            w186=> c0_n43_w186, 
            w187=> c0_n43_w187, 
            w188=> c0_n43_w188, 
            w189=> c0_n43_w189, 
            w190=> c0_n43_w190, 
            w191=> c0_n43_w191, 
            w192=> c0_n43_w192, 
            w193=> c0_n43_w193, 
            w194=> c0_n43_w194, 
            w195=> c0_n43_w195, 
            w196=> c0_n43_w196, 
            w197=> c0_n43_w197, 
            w198=> c0_n43_w198, 
            w199=> c0_n43_w199, 
            w200=> c0_n43_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n43_y
   );           
            
neuron_inst_44: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n44_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n44_w1, 
            w2=> c0_n44_w2, 
            w3=> c0_n44_w3, 
            w4=> c0_n44_w4, 
            w5=> c0_n44_w5, 
            w6=> c0_n44_w6, 
            w7=> c0_n44_w7, 
            w8=> c0_n44_w8, 
            w9=> c0_n44_w9, 
            w10=> c0_n44_w10, 
            w11=> c0_n44_w11, 
            w12=> c0_n44_w12, 
            w13=> c0_n44_w13, 
            w14=> c0_n44_w14, 
            w15=> c0_n44_w15, 
            w16=> c0_n44_w16, 
            w17=> c0_n44_w17, 
            w18=> c0_n44_w18, 
            w19=> c0_n44_w19, 
            w20=> c0_n44_w20, 
            w21=> c0_n44_w21, 
            w22=> c0_n44_w22, 
            w23=> c0_n44_w23, 
            w24=> c0_n44_w24, 
            w25=> c0_n44_w25, 
            w26=> c0_n44_w26, 
            w27=> c0_n44_w27, 
            w28=> c0_n44_w28, 
            w29=> c0_n44_w29, 
            w30=> c0_n44_w30, 
            w31=> c0_n44_w31, 
            w32=> c0_n44_w32, 
            w33=> c0_n44_w33, 
            w34=> c0_n44_w34, 
            w35=> c0_n44_w35, 
            w36=> c0_n44_w36, 
            w37=> c0_n44_w37, 
            w38=> c0_n44_w38, 
            w39=> c0_n44_w39, 
            w40=> c0_n44_w40, 
            w41=> c0_n44_w41, 
            w42=> c0_n44_w42, 
            w43=> c0_n44_w43, 
            w44=> c0_n44_w44, 
            w45=> c0_n44_w45, 
            w46=> c0_n44_w46, 
            w47=> c0_n44_w47, 
            w48=> c0_n44_w48, 
            w49=> c0_n44_w49, 
            w50=> c0_n44_w50, 
            w51=> c0_n44_w51, 
            w52=> c0_n44_w52, 
            w53=> c0_n44_w53, 
            w54=> c0_n44_w54, 
            w55=> c0_n44_w55, 
            w56=> c0_n44_w56, 
            w57=> c0_n44_w57, 
            w58=> c0_n44_w58, 
            w59=> c0_n44_w59, 
            w60=> c0_n44_w60, 
            w61=> c0_n44_w61, 
            w62=> c0_n44_w62, 
            w63=> c0_n44_w63, 
            w64=> c0_n44_w64, 
            w65=> c0_n44_w65, 
            w66=> c0_n44_w66, 
            w67=> c0_n44_w67, 
            w68=> c0_n44_w68, 
            w69=> c0_n44_w69, 
            w70=> c0_n44_w70, 
            w71=> c0_n44_w71, 
            w72=> c0_n44_w72, 
            w73=> c0_n44_w73, 
            w74=> c0_n44_w74, 
            w75=> c0_n44_w75, 
            w76=> c0_n44_w76, 
            w77=> c0_n44_w77, 
            w78=> c0_n44_w78, 
            w79=> c0_n44_w79, 
            w80=> c0_n44_w80, 
            w81=> c0_n44_w81, 
            w82=> c0_n44_w82, 
            w83=> c0_n44_w83, 
            w84=> c0_n44_w84, 
            w85=> c0_n44_w85, 
            w86=> c0_n44_w86, 
            w87=> c0_n44_w87, 
            w88=> c0_n44_w88, 
            w89=> c0_n44_w89, 
            w90=> c0_n44_w90, 
            w91=> c0_n44_w91, 
            w92=> c0_n44_w92, 
            w93=> c0_n44_w93, 
            w94=> c0_n44_w94, 
            w95=> c0_n44_w95, 
            w96=> c0_n44_w96, 
            w97=> c0_n44_w97, 
            w98=> c0_n44_w98, 
            w99=> c0_n44_w99, 
            w100=> c0_n44_w100, 
            w101=> c0_n44_w101, 
            w102=> c0_n44_w102, 
            w103=> c0_n44_w103, 
            w104=> c0_n44_w104, 
            w105=> c0_n44_w105, 
            w106=> c0_n44_w106, 
            w107=> c0_n44_w107, 
            w108=> c0_n44_w108, 
            w109=> c0_n44_w109, 
            w110=> c0_n44_w110, 
            w111=> c0_n44_w111, 
            w112=> c0_n44_w112, 
            w113=> c0_n44_w113, 
            w114=> c0_n44_w114, 
            w115=> c0_n44_w115, 
            w116=> c0_n44_w116, 
            w117=> c0_n44_w117, 
            w118=> c0_n44_w118, 
            w119=> c0_n44_w119, 
            w120=> c0_n44_w120, 
            w121=> c0_n44_w121, 
            w122=> c0_n44_w122, 
            w123=> c0_n44_w123, 
            w124=> c0_n44_w124, 
            w125=> c0_n44_w125, 
            w126=> c0_n44_w126, 
            w127=> c0_n44_w127, 
            w128=> c0_n44_w128, 
            w129=> c0_n44_w129, 
            w130=> c0_n44_w130, 
            w131=> c0_n44_w131, 
            w132=> c0_n44_w132, 
            w133=> c0_n44_w133, 
            w134=> c0_n44_w134, 
            w135=> c0_n44_w135, 
            w136=> c0_n44_w136, 
            w137=> c0_n44_w137, 
            w138=> c0_n44_w138, 
            w139=> c0_n44_w139, 
            w140=> c0_n44_w140, 
            w141=> c0_n44_w141, 
            w142=> c0_n44_w142, 
            w143=> c0_n44_w143, 
            w144=> c0_n44_w144, 
            w145=> c0_n44_w145, 
            w146=> c0_n44_w146, 
            w147=> c0_n44_w147, 
            w148=> c0_n44_w148, 
            w149=> c0_n44_w149, 
            w150=> c0_n44_w150, 
            w151=> c0_n44_w151, 
            w152=> c0_n44_w152, 
            w153=> c0_n44_w153, 
            w154=> c0_n44_w154, 
            w155=> c0_n44_w155, 
            w156=> c0_n44_w156, 
            w157=> c0_n44_w157, 
            w158=> c0_n44_w158, 
            w159=> c0_n44_w159, 
            w160=> c0_n44_w160, 
            w161=> c0_n44_w161, 
            w162=> c0_n44_w162, 
            w163=> c0_n44_w163, 
            w164=> c0_n44_w164, 
            w165=> c0_n44_w165, 
            w166=> c0_n44_w166, 
            w167=> c0_n44_w167, 
            w168=> c0_n44_w168, 
            w169=> c0_n44_w169, 
            w170=> c0_n44_w170, 
            w171=> c0_n44_w171, 
            w172=> c0_n44_w172, 
            w173=> c0_n44_w173, 
            w174=> c0_n44_w174, 
            w175=> c0_n44_w175, 
            w176=> c0_n44_w176, 
            w177=> c0_n44_w177, 
            w178=> c0_n44_w178, 
            w179=> c0_n44_w179, 
            w180=> c0_n44_w180, 
            w181=> c0_n44_w181, 
            w182=> c0_n44_w182, 
            w183=> c0_n44_w183, 
            w184=> c0_n44_w184, 
            w185=> c0_n44_w185, 
            w186=> c0_n44_w186, 
            w187=> c0_n44_w187, 
            w188=> c0_n44_w188, 
            w189=> c0_n44_w189, 
            w190=> c0_n44_w190, 
            w191=> c0_n44_w191, 
            w192=> c0_n44_w192, 
            w193=> c0_n44_w193, 
            w194=> c0_n44_w194, 
            w195=> c0_n44_w195, 
            w196=> c0_n44_w196, 
            w197=> c0_n44_w197, 
            w198=> c0_n44_w198, 
            w199=> c0_n44_w199, 
            w200=> c0_n44_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n44_y
   );           
            
neuron_inst_45: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n45_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n45_w1, 
            w2=> c0_n45_w2, 
            w3=> c0_n45_w3, 
            w4=> c0_n45_w4, 
            w5=> c0_n45_w5, 
            w6=> c0_n45_w6, 
            w7=> c0_n45_w7, 
            w8=> c0_n45_w8, 
            w9=> c0_n45_w9, 
            w10=> c0_n45_w10, 
            w11=> c0_n45_w11, 
            w12=> c0_n45_w12, 
            w13=> c0_n45_w13, 
            w14=> c0_n45_w14, 
            w15=> c0_n45_w15, 
            w16=> c0_n45_w16, 
            w17=> c0_n45_w17, 
            w18=> c0_n45_w18, 
            w19=> c0_n45_w19, 
            w20=> c0_n45_w20, 
            w21=> c0_n45_w21, 
            w22=> c0_n45_w22, 
            w23=> c0_n45_w23, 
            w24=> c0_n45_w24, 
            w25=> c0_n45_w25, 
            w26=> c0_n45_w26, 
            w27=> c0_n45_w27, 
            w28=> c0_n45_w28, 
            w29=> c0_n45_w29, 
            w30=> c0_n45_w30, 
            w31=> c0_n45_w31, 
            w32=> c0_n45_w32, 
            w33=> c0_n45_w33, 
            w34=> c0_n45_w34, 
            w35=> c0_n45_w35, 
            w36=> c0_n45_w36, 
            w37=> c0_n45_w37, 
            w38=> c0_n45_w38, 
            w39=> c0_n45_w39, 
            w40=> c0_n45_w40, 
            w41=> c0_n45_w41, 
            w42=> c0_n45_w42, 
            w43=> c0_n45_w43, 
            w44=> c0_n45_w44, 
            w45=> c0_n45_w45, 
            w46=> c0_n45_w46, 
            w47=> c0_n45_w47, 
            w48=> c0_n45_w48, 
            w49=> c0_n45_w49, 
            w50=> c0_n45_w50, 
            w51=> c0_n45_w51, 
            w52=> c0_n45_w52, 
            w53=> c0_n45_w53, 
            w54=> c0_n45_w54, 
            w55=> c0_n45_w55, 
            w56=> c0_n45_w56, 
            w57=> c0_n45_w57, 
            w58=> c0_n45_w58, 
            w59=> c0_n45_w59, 
            w60=> c0_n45_w60, 
            w61=> c0_n45_w61, 
            w62=> c0_n45_w62, 
            w63=> c0_n45_w63, 
            w64=> c0_n45_w64, 
            w65=> c0_n45_w65, 
            w66=> c0_n45_w66, 
            w67=> c0_n45_w67, 
            w68=> c0_n45_w68, 
            w69=> c0_n45_w69, 
            w70=> c0_n45_w70, 
            w71=> c0_n45_w71, 
            w72=> c0_n45_w72, 
            w73=> c0_n45_w73, 
            w74=> c0_n45_w74, 
            w75=> c0_n45_w75, 
            w76=> c0_n45_w76, 
            w77=> c0_n45_w77, 
            w78=> c0_n45_w78, 
            w79=> c0_n45_w79, 
            w80=> c0_n45_w80, 
            w81=> c0_n45_w81, 
            w82=> c0_n45_w82, 
            w83=> c0_n45_w83, 
            w84=> c0_n45_w84, 
            w85=> c0_n45_w85, 
            w86=> c0_n45_w86, 
            w87=> c0_n45_w87, 
            w88=> c0_n45_w88, 
            w89=> c0_n45_w89, 
            w90=> c0_n45_w90, 
            w91=> c0_n45_w91, 
            w92=> c0_n45_w92, 
            w93=> c0_n45_w93, 
            w94=> c0_n45_w94, 
            w95=> c0_n45_w95, 
            w96=> c0_n45_w96, 
            w97=> c0_n45_w97, 
            w98=> c0_n45_w98, 
            w99=> c0_n45_w99, 
            w100=> c0_n45_w100, 
            w101=> c0_n45_w101, 
            w102=> c0_n45_w102, 
            w103=> c0_n45_w103, 
            w104=> c0_n45_w104, 
            w105=> c0_n45_w105, 
            w106=> c0_n45_w106, 
            w107=> c0_n45_w107, 
            w108=> c0_n45_w108, 
            w109=> c0_n45_w109, 
            w110=> c0_n45_w110, 
            w111=> c0_n45_w111, 
            w112=> c0_n45_w112, 
            w113=> c0_n45_w113, 
            w114=> c0_n45_w114, 
            w115=> c0_n45_w115, 
            w116=> c0_n45_w116, 
            w117=> c0_n45_w117, 
            w118=> c0_n45_w118, 
            w119=> c0_n45_w119, 
            w120=> c0_n45_w120, 
            w121=> c0_n45_w121, 
            w122=> c0_n45_w122, 
            w123=> c0_n45_w123, 
            w124=> c0_n45_w124, 
            w125=> c0_n45_w125, 
            w126=> c0_n45_w126, 
            w127=> c0_n45_w127, 
            w128=> c0_n45_w128, 
            w129=> c0_n45_w129, 
            w130=> c0_n45_w130, 
            w131=> c0_n45_w131, 
            w132=> c0_n45_w132, 
            w133=> c0_n45_w133, 
            w134=> c0_n45_w134, 
            w135=> c0_n45_w135, 
            w136=> c0_n45_w136, 
            w137=> c0_n45_w137, 
            w138=> c0_n45_w138, 
            w139=> c0_n45_w139, 
            w140=> c0_n45_w140, 
            w141=> c0_n45_w141, 
            w142=> c0_n45_w142, 
            w143=> c0_n45_w143, 
            w144=> c0_n45_w144, 
            w145=> c0_n45_w145, 
            w146=> c0_n45_w146, 
            w147=> c0_n45_w147, 
            w148=> c0_n45_w148, 
            w149=> c0_n45_w149, 
            w150=> c0_n45_w150, 
            w151=> c0_n45_w151, 
            w152=> c0_n45_w152, 
            w153=> c0_n45_w153, 
            w154=> c0_n45_w154, 
            w155=> c0_n45_w155, 
            w156=> c0_n45_w156, 
            w157=> c0_n45_w157, 
            w158=> c0_n45_w158, 
            w159=> c0_n45_w159, 
            w160=> c0_n45_w160, 
            w161=> c0_n45_w161, 
            w162=> c0_n45_w162, 
            w163=> c0_n45_w163, 
            w164=> c0_n45_w164, 
            w165=> c0_n45_w165, 
            w166=> c0_n45_w166, 
            w167=> c0_n45_w167, 
            w168=> c0_n45_w168, 
            w169=> c0_n45_w169, 
            w170=> c0_n45_w170, 
            w171=> c0_n45_w171, 
            w172=> c0_n45_w172, 
            w173=> c0_n45_w173, 
            w174=> c0_n45_w174, 
            w175=> c0_n45_w175, 
            w176=> c0_n45_w176, 
            w177=> c0_n45_w177, 
            w178=> c0_n45_w178, 
            w179=> c0_n45_w179, 
            w180=> c0_n45_w180, 
            w181=> c0_n45_w181, 
            w182=> c0_n45_w182, 
            w183=> c0_n45_w183, 
            w184=> c0_n45_w184, 
            w185=> c0_n45_w185, 
            w186=> c0_n45_w186, 
            w187=> c0_n45_w187, 
            w188=> c0_n45_w188, 
            w189=> c0_n45_w189, 
            w190=> c0_n45_w190, 
            w191=> c0_n45_w191, 
            w192=> c0_n45_w192, 
            w193=> c0_n45_w193, 
            w194=> c0_n45_w194, 
            w195=> c0_n45_w195, 
            w196=> c0_n45_w196, 
            w197=> c0_n45_w197, 
            w198=> c0_n45_w198, 
            w199=> c0_n45_w199, 
            w200=> c0_n45_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n45_y
   );           
            
neuron_inst_46: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n46_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n46_w1, 
            w2=> c0_n46_w2, 
            w3=> c0_n46_w3, 
            w4=> c0_n46_w4, 
            w5=> c0_n46_w5, 
            w6=> c0_n46_w6, 
            w7=> c0_n46_w7, 
            w8=> c0_n46_w8, 
            w9=> c0_n46_w9, 
            w10=> c0_n46_w10, 
            w11=> c0_n46_w11, 
            w12=> c0_n46_w12, 
            w13=> c0_n46_w13, 
            w14=> c0_n46_w14, 
            w15=> c0_n46_w15, 
            w16=> c0_n46_w16, 
            w17=> c0_n46_w17, 
            w18=> c0_n46_w18, 
            w19=> c0_n46_w19, 
            w20=> c0_n46_w20, 
            w21=> c0_n46_w21, 
            w22=> c0_n46_w22, 
            w23=> c0_n46_w23, 
            w24=> c0_n46_w24, 
            w25=> c0_n46_w25, 
            w26=> c0_n46_w26, 
            w27=> c0_n46_w27, 
            w28=> c0_n46_w28, 
            w29=> c0_n46_w29, 
            w30=> c0_n46_w30, 
            w31=> c0_n46_w31, 
            w32=> c0_n46_w32, 
            w33=> c0_n46_w33, 
            w34=> c0_n46_w34, 
            w35=> c0_n46_w35, 
            w36=> c0_n46_w36, 
            w37=> c0_n46_w37, 
            w38=> c0_n46_w38, 
            w39=> c0_n46_w39, 
            w40=> c0_n46_w40, 
            w41=> c0_n46_w41, 
            w42=> c0_n46_w42, 
            w43=> c0_n46_w43, 
            w44=> c0_n46_w44, 
            w45=> c0_n46_w45, 
            w46=> c0_n46_w46, 
            w47=> c0_n46_w47, 
            w48=> c0_n46_w48, 
            w49=> c0_n46_w49, 
            w50=> c0_n46_w50, 
            w51=> c0_n46_w51, 
            w52=> c0_n46_w52, 
            w53=> c0_n46_w53, 
            w54=> c0_n46_w54, 
            w55=> c0_n46_w55, 
            w56=> c0_n46_w56, 
            w57=> c0_n46_w57, 
            w58=> c0_n46_w58, 
            w59=> c0_n46_w59, 
            w60=> c0_n46_w60, 
            w61=> c0_n46_w61, 
            w62=> c0_n46_w62, 
            w63=> c0_n46_w63, 
            w64=> c0_n46_w64, 
            w65=> c0_n46_w65, 
            w66=> c0_n46_w66, 
            w67=> c0_n46_w67, 
            w68=> c0_n46_w68, 
            w69=> c0_n46_w69, 
            w70=> c0_n46_w70, 
            w71=> c0_n46_w71, 
            w72=> c0_n46_w72, 
            w73=> c0_n46_w73, 
            w74=> c0_n46_w74, 
            w75=> c0_n46_w75, 
            w76=> c0_n46_w76, 
            w77=> c0_n46_w77, 
            w78=> c0_n46_w78, 
            w79=> c0_n46_w79, 
            w80=> c0_n46_w80, 
            w81=> c0_n46_w81, 
            w82=> c0_n46_w82, 
            w83=> c0_n46_w83, 
            w84=> c0_n46_w84, 
            w85=> c0_n46_w85, 
            w86=> c0_n46_w86, 
            w87=> c0_n46_w87, 
            w88=> c0_n46_w88, 
            w89=> c0_n46_w89, 
            w90=> c0_n46_w90, 
            w91=> c0_n46_w91, 
            w92=> c0_n46_w92, 
            w93=> c0_n46_w93, 
            w94=> c0_n46_w94, 
            w95=> c0_n46_w95, 
            w96=> c0_n46_w96, 
            w97=> c0_n46_w97, 
            w98=> c0_n46_w98, 
            w99=> c0_n46_w99, 
            w100=> c0_n46_w100, 
            w101=> c0_n46_w101, 
            w102=> c0_n46_w102, 
            w103=> c0_n46_w103, 
            w104=> c0_n46_w104, 
            w105=> c0_n46_w105, 
            w106=> c0_n46_w106, 
            w107=> c0_n46_w107, 
            w108=> c0_n46_w108, 
            w109=> c0_n46_w109, 
            w110=> c0_n46_w110, 
            w111=> c0_n46_w111, 
            w112=> c0_n46_w112, 
            w113=> c0_n46_w113, 
            w114=> c0_n46_w114, 
            w115=> c0_n46_w115, 
            w116=> c0_n46_w116, 
            w117=> c0_n46_w117, 
            w118=> c0_n46_w118, 
            w119=> c0_n46_w119, 
            w120=> c0_n46_w120, 
            w121=> c0_n46_w121, 
            w122=> c0_n46_w122, 
            w123=> c0_n46_w123, 
            w124=> c0_n46_w124, 
            w125=> c0_n46_w125, 
            w126=> c0_n46_w126, 
            w127=> c0_n46_w127, 
            w128=> c0_n46_w128, 
            w129=> c0_n46_w129, 
            w130=> c0_n46_w130, 
            w131=> c0_n46_w131, 
            w132=> c0_n46_w132, 
            w133=> c0_n46_w133, 
            w134=> c0_n46_w134, 
            w135=> c0_n46_w135, 
            w136=> c0_n46_w136, 
            w137=> c0_n46_w137, 
            w138=> c0_n46_w138, 
            w139=> c0_n46_w139, 
            w140=> c0_n46_w140, 
            w141=> c0_n46_w141, 
            w142=> c0_n46_w142, 
            w143=> c0_n46_w143, 
            w144=> c0_n46_w144, 
            w145=> c0_n46_w145, 
            w146=> c0_n46_w146, 
            w147=> c0_n46_w147, 
            w148=> c0_n46_w148, 
            w149=> c0_n46_w149, 
            w150=> c0_n46_w150, 
            w151=> c0_n46_w151, 
            w152=> c0_n46_w152, 
            w153=> c0_n46_w153, 
            w154=> c0_n46_w154, 
            w155=> c0_n46_w155, 
            w156=> c0_n46_w156, 
            w157=> c0_n46_w157, 
            w158=> c0_n46_w158, 
            w159=> c0_n46_w159, 
            w160=> c0_n46_w160, 
            w161=> c0_n46_w161, 
            w162=> c0_n46_w162, 
            w163=> c0_n46_w163, 
            w164=> c0_n46_w164, 
            w165=> c0_n46_w165, 
            w166=> c0_n46_w166, 
            w167=> c0_n46_w167, 
            w168=> c0_n46_w168, 
            w169=> c0_n46_w169, 
            w170=> c0_n46_w170, 
            w171=> c0_n46_w171, 
            w172=> c0_n46_w172, 
            w173=> c0_n46_w173, 
            w174=> c0_n46_w174, 
            w175=> c0_n46_w175, 
            w176=> c0_n46_w176, 
            w177=> c0_n46_w177, 
            w178=> c0_n46_w178, 
            w179=> c0_n46_w179, 
            w180=> c0_n46_w180, 
            w181=> c0_n46_w181, 
            w182=> c0_n46_w182, 
            w183=> c0_n46_w183, 
            w184=> c0_n46_w184, 
            w185=> c0_n46_w185, 
            w186=> c0_n46_w186, 
            w187=> c0_n46_w187, 
            w188=> c0_n46_w188, 
            w189=> c0_n46_w189, 
            w190=> c0_n46_w190, 
            w191=> c0_n46_w191, 
            w192=> c0_n46_w192, 
            w193=> c0_n46_w193, 
            w194=> c0_n46_w194, 
            w195=> c0_n46_w195, 
            w196=> c0_n46_w196, 
            w197=> c0_n46_w197, 
            w198=> c0_n46_w198, 
            w199=> c0_n46_w199, 
            w200=> c0_n46_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n46_y
   );           
            
neuron_inst_47: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n47_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n47_w1, 
            w2=> c0_n47_w2, 
            w3=> c0_n47_w3, 
            w4=> c0_n47_w4, 
            w5=> c0_n47_w5, 
            w6=> c0_n47_w6, 
            w7=> c0_n47_w7, 
            w8=> c0_n47_w8, 
            w9=> c0_n47_w9, 
            w10=> c0_n47_w10, 
            w11=> c0_n47_w11, 
            w12=> c0_n47_w12, 
            w13=> c0_n47_w13, 
            w14=> c0_n47_w14, 
            w15=> c0_n47_w15, 
            w16=> c0_n47_w16, 
            w17=> c0_n47_w17, 
            w18=> c0_n47_w18, 
            w19=> c0_n47_w19, 
            w20=> c0_n47_w20, 
            w21=> c0_n47_w21, 
            w22=> c0_n47_w22, 
            w23=> c0_n47_w23, 
            w24=> c0_n47_w24, 
            w25=> c0_n47_w25, 
            w26=> c0_n47_w26, 
            w27=> c0_n47_w27, 
            w28=> c0_n47_w28, 
            w29=> c0_n47_w29, 
            w30=> c0_n47_w30, 
            w31=> c0_n47_w31, 
            w32=> c0_n47_w32, 
            w33=> c0_n47_w33, 
            w34=> c0_n47_w34, 
            w35=> c0_n47_w35, 
            w36=> c0_n47_w36, 
            w37=> c0_n47_w37, 
            w38=> c0_n47_w38, 
            w39=> c0_n47_w39, 
            w40=> c0_n47_w40, 
            w41=> c0_n47_w41, 
            w42=> c0_n47_w42, 
            w43=> c0_n47_w43, 
            w44=> c0_n47_w44, 
            w45=> c0_n47_w45, 
            w46=> c0_n47_w46, 
            w47=> c0_n47_w47, 
            w48=> c0_n47_w48, 
            w49=> c0_n47_w49, 
            w50=> c0_n47_w50, 
            w51=> c0_n47_w51, 
            w52=> c0_n47_w52, 
            w53=> c0_n47_w53, 
            w54=> c0_n47_w54, 
            w55=> c0_n47_w55, 
            w56=> c0_n47_w56, 
            w57=> c0_n47_w57, 
            w58=> c0_n47_w58, 
            w59=> c0_n47_w59, 
            w60=> c0_n47_w60, 
            w61=> c0_n47_w61, 
            w62=> c0_n47_w62, 
            w63=> c0_n47_w63, 
            w64=> c0_n47_w64, 
            w65=> c0_n47_w65, 
            w66=> c0_n47_w66, 
            w67=> c0_n47_w67, 
            w68=> c0_n47_w68, 
            w69=> c0_n47_w69, 
            w70=> c0_n47_w70, 
            w71=> c0_n47_w71, 
            w72=> c0_n47_w72, 
            w73=> c0_n47_w73, 
            w74=> c0_n47_w74, 
            w75=> c0_n47_w75, 
            w76=> c0_n47_w76, 
            w77=> c0_n47_w77, 
            w78=> c0_n47_w78, 
            w79=> c0_n47_w79, 
            w80=> c0_n47_w80, 
            w81=> c0_n47_w81, 
            w82=> c0_n47_w82, 
            w83=> c0_n47_w83, 
            w84=> c0_n47_w84, 
            w85=> c0_n47_w85, 
            w86=> c0_n47_w86, 
            w87=> c0_n47_w87, 
            w88=> c0_n47_w88, 
            w89=> c0_n47_w89, 
            w90=> c0_n47_w90, 
            w91=> c0_n47_w91, 
            w92=> c0_n47_w92, 
            w93=> c0_n47_w93, 
            w94=> c0_n47_w94, 
            w95=> c0_n47_w95, 
            w96=> c0_n47_w96, 
            w97=> c0_n47_w97, 
            w98=> c0_n47_w98, 
            w99=> c0_n47_w99, 
            w100=> c0_n47_w100, 
            w101=> c0_n47_w101, 
            w102=> c0_n47_w102, 
            w103=> c0_n47_w103, 
            w104=> c0_n47_w104, 
            w105=> c0_n47_w105, 
            w106=> c0_n47_w106, 
            w107=> c0_n47_w107, 
            w108=> c0_n47_w108, 
            w109=> c0_n47_w109, 
            w110=> c0_n47_w110, 
            w111=> c0_n47_w111, 
            w112=> c0_n47_w112, 
            w113=> c0_n47_w113, 
            w114=> c0_n47_w114, 
            w115=> c0_n47_w115, 
            w116=> c0_n47_w116, 
            w117=> c0_n47_w117, 
            w118=> c0_n47_w118, 
            w119=> c0_n47_w119, 
            w120=> c0_n47_w120, 
            w121=> c0_n47_w121, 
            w122=> c0_n47_w122, 
            w123=> c0_n47_w123, 
            w124=> c0_n47_w124, 
            w125=> c0_n47_w125, 
            w126=> c0_n47_w126, 
            w127=> c0_n47_w127, 
            w128=> c0_n47_w128, 
            w129=> c0_n47_w129, 
            w130=> c0_n47_w130, 
            w131=> c0_n47_w131, 
            w132=> c0_n47_w132, 
            w133=> c0_n47_w133, 
            w134=> c0_n47_w134, 
            w135=> c0_n47_w135, 
            w136=> c0_n47_w136, 
            w137=> c0_n47_w137, 
            w138=> c0_n47_w138, 
            w139=> c0_n47_w139, 
            w140=> c0_n47_w140, 
            w141=> c0_n47_w141, 
            w142=> c0_n47_w142, 
            w143=> c0_n47_w143, 
            w144=> c0_n47_w144, 
            w145=> c0_n47_w145, 
            w146=> c0_n47_w146, 
            w147=> c0_n47_w147, 
            w148=> c0_n47_w148, 
            w149=> c0_n47_w149, 
            w150=> c0_n47_w150, 
            w151=> c0_n47_w151, 
            w152=> c0_n47_w152, 
            w153=> c0_n47_w153, 
            w154=> c0_n47_w154, 
            w155=> c0_n47_w155, 
            w156=> c0_n47_w156, 
            w157=> c0_n47_w157, 
            w158=> c0_n47_w158, 
            w159=> c0_n47_w159, 
            w160=> c0_n47_w160, 
            w161=> c0_n47_w161, 
            w162=> c0_n47_w162, 
            w163=> c0_n47_w163, 
            w164=> c0_n47_w164, 
            w165=> c0_n47_w165, 
            w166=> c0_n47_w166, 
            w167=> c0_n47_w167, 
            w168=> c0_n47_w168, 
            w169=> c0_n47_w169, 
            w170=> c0_n47_w170, 
            w171=> c0_n47_w171, 
            w172=> c0_n47_w172, 
            w173=> c0_n47_w173, 
            w174=> c0_n47_w174, 
            w175=> c0_n47_w175, 
            w176=> c0_n47_w176, 
            w177=> c0_n47_w177, 
            w178=> c0_n47_w178, 
            w179=> c0_n47_w179, 
            w180=> c0_n47_w180, 
            w181=> c0_n47_w181, 
            w182=> c0_n47_w182, 
            w183=> c0_n47_w183, 
            w184=> c0_n47_w184, 
            w185=> c0_n47_w185, 
            w186=> c0_n47_w186, 
            w187=> c0_n47_w187, 
            w188=> c0_n47_w188, 
            w189=> c0_n47_w189, 
            w190=> c0_n47_w190, 
            w191=> c0_n47_w191, 
            w192=> c0_n47_w192, 
            w193=> c0_n47_w193, 
            w194=> c0_n47_w194, 
            w195=> c0_n47_w195, 
            w196=> c0_n47_w196, 
            w197=> c0_n47_w197, 
            w198=> c0_n47_w198, 
            w199=> c0_n47_w199, 
            w200=> c0_n47_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n47_y
   );           
            
neuron_inst_48: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n48_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n48_w1, 
            w2=> c0_n48_w2, 
            w3=> c0_n48_w3, 
            w4=> c0_n48_w4, 
            w5=> c0_n48_w5, 
            w6=> c0_n48_w6, 
            w7=> c0_n48_w7, 
            w8=> c0_n48_w8, 
            w9=> c0_n48_w9, 
            w10=> c0_n48_w10, 
            w11=> c0_n48_w11, 
            w12=> c0_n48_w12, 
            w13=> c0_n48_w13, 
            w14=> c0_n48_w14, 
            w15=> c0_n48_w15, 
            w16=> c0_n48_w16, 
            w17=> c0_n48_w17, 
            w18=> c0_n48_w18, 
            w19=> c0_n48_w19, 
            w20=> c0_n48_w20, 
            w21=> c0_n48_w21, 
            w22=> c0_n48_w22, 
            w23=> c0_n48_w23, 
            w24=> c0_n48_w24, 
            w25=> c0_n48_w25, 
            w26=> c0_n48_w26, 
            w27=> c0_n48_w27, 
            w28=> c0_n48_w28, 
            w29=> c0_n48_w29, 
            w30=> c0_n48_w30, 
            w31=> c0_n48_w31, 
            w32=> c0_n48_w32, 
            w33=> c0_n48_w33, 
            w34=> c0_n48_w34, 
            w35=> c0_n48_w35, 
            w36=> c0_n48_w36, 
            w37=> c0_n48_w37, 
            w38=> c0_n48_w38, 
            w39=> c0_n48_w39, 
            w40=> c0_n48_w40, 
            w41=> c0_n48_w41, 
            w42=> c0_n48_w42, 
            w43=> c0_n48_w43, 
            w44=> c0_n48_w44, 
            w45=> c0_n48_w45, 
            w46=> c0_n48_w46, 
            w47=> c0_n48_w47, 
            w48=> c0_n48_w48, 
            w49=> c0_n48_w49, 
            w50=> c0_n48_w50, 
            w51=> c0_n48_w51, 
            w52=> c0_n48_w52, 
            w53=> c0_n48_w53, 
            w54=> c0_n48_w54, 
            w55=> c0_n48_w55, 
            w56=> c0_n48_w56, 
            w57=> c0_n48_w57, 
            w58=> c0_n48_w58, 
            w59=> c0_n48_w59, 
            w60=> c0_n48_w60, 
            w61=> c0_n48_w61, 
            w62=> c0_n48_w62, 
            w63=> c0_n48_w63, 
            w64=> c0_n48_w64, 
            w65=> c0_n48_w65, 
            w66=> c0_n48_w66, 
            w67=> c0_n48_w67, 
            w68=> c0_n48_w68, 
            w69=> c0_n48_w69, 
            w70=> c0_n48_w70, 
            w71=> c0_n48_w71, 
            w72=> c0_n48_w72, 
            w73=> c0_n48_w73, 
            w74=> c0_n48_w74, 
            w75=> c0_n48_w75, 
            w76=> c0_n48_w76, 
            w77=> c0_n48_w77, 
            w78=> c0_n48_w78, 
            w79=> c0_n48_w79, 
            w80=> c0_n48_w80, 
            w81=> c0_n48_w81, 
            w82=> c0_n48_w82, 
            w83=> c0_n48_w83, 
            w84=> c0_n48_w84, 
            w85=> c0_n48_w85, 
            w86=> c0_n48_w86, 
            w87=> c0_n48_w87, 
            w88=> c0_n48_w88, 
            w89=> c0_n48_w89, 
            w90=> c0_n48_w90, 
            w91=> c0_n48_w91, 
            w92=> c0_n48_w92, 
            w93=> c0_n48_w93, 
            w94=> c0_n48_w94, 
            w95=> c0_n48_w95, 
            w96=> c0_n48_w96, 
            w97=> c0_n48_w97, 
            w98=> c0_n48_w98, 
            w99=> c0_n48_w99, 
            w100=> c0_n48_w100, 
            w101=> c0_n48_w101, 
            w102=> c0_n48_w102, 
            w103=> c0_n48_w103, 
            w104=> c0_n48_w104, 
            w105=> c0_n48_w105, 
            w106=> c0_n48_w106, 
            w107=> c0_n48_w107, 
            w108=> c0_n48_w108, 
            w109=> c0_n48_w109, 
            w110=> c0_n48_w110, 
            w111=> c0_n48_w111, 
            w112=> c0_n48_w112, 
            w113=> c0_n48_w113, 
            w114=> c0_n48_w114, 
            w115=> c0_n48_w115, 
            w116=> c0_n48_w116, 
            w117=> c0_n48_w117, 
            w118=> c0_n48_w118, 
            w119=> c0_n48_w119, 
            w120=> c0_n48_w120, 
            w121=> c0_n48_w121, 
            w122=> c0_n48_w122, 
            w123=> c0_n48_w123, 
            w124=> c0_n48_w124, 
            w125=> c0_n48_w125, 
            w126=> c0_n48_w126, 
            w127=> c0_n48_w127, 
            w128=> c0_n48_w128, 
            w129=> c0_n48_w129, 
            w130=> c0_n48_w130, 
            w131=> c0_n48_w131, 
            w132=> c0_n48_w132, 
            w133=> c0_n48_w133, 
            w134=> c0_n48_w134, 
            w135=> c0_n48_w135, 
            w136=> c0_n48_w136, 
            w137=> c0_n48_w137, 
            w138=> c0_n48_w138, 
            w139=> c0_n48_w139, 
            w140=> c0_n48_w140, 
            w141=> c0_n48_w141, 
            w142=> c0_n48_w142, 
            w143=> c0_n48_w143, 
            w144=> c0_n48_w144, 
            w145=> c0_n48_w145, 
            w146=> c0_n48_w146, 
            w147=> c0_n48_w147, 
            w148=> c0_n48_w148, 
            w149=> c0_n48_w149, 
            w150=> c0_n48_w150, 
            w151=> c0_n48_w151, 
            w152=> c0_n48_w152, 
            w153=> c0_n48_w153, 
            w154=> c0_n48_w154, 
            w155=> c0_n48_w155, 
            w156=> c0_n48_w156, 
            w157=> c0_n48_w157, 
            w158=> c0_n48_w158, 
            w159=> c0_n48_w159, 
            w160=> c0_n48_w160, 
            w161=> c0_n48_w161, 
            w162=> c0_n48_w162, 
            w163=> c0_n48_w163, 
            w164=> c0_n48_w164, 
            w165=> c0_n48_w165, 
            w166=> c0_n48_w166, 
            w167=> c0_n48_w167, 
            w168=> c0_n48_w168, 
            w169=> c0_n48_w169, 
            w170=> c0_n48_w170, 
            w171=> c0_n48_w171, 
            w172=> c0_n48_w172, 
            w173=> c0_n48_w173, 
            w174=> c0_n48_w174, 
            w175=> c0_n48_w175, 
            w176=> c0_n48_w176, 
            w177=> c0_n48_w177, 
            w178=> c0_n48_w178, 
            w179=> c0_n48_w179, 
            w180=> c0_n48_w180, 
            w181=> c0_n48_w181, 
            w182=> c0_n48_w182, 
            w183=> c0_n48_w183, 
            w184=> c0_n48_w184, 
            w185=> c0_n48_w185, 
            w186=> c0_n48_w186, 
            w187=> c0_n48_w187, 
            w188=> c0_n48_w188, 
            w189=> c0_n48_w189, 
            w190=> c0_n48_w190, 
            w191=> c0_n48_w191, 
            w192=> c0_n48_w192, 
            w193=> c0_n48_w193, 
            w194=> c0_n48_w194, 
            w195=> c0_n48_w195, 
            w196=> c0_n48_w196, 
            w197=> c0_n48_w197, 
            w198=> c0_n48_w198, 
            w199=> c0_n48_w199, 
            w200=> c0_n48_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n48_y
   );           
            
neuron_inst_49: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n49_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n49_w1, 
            w2=> c0_n49_w2, 
            w3=> c0_n49_w3, 
            w4=> c0_n49_w4, 
            w5=> c0_n49_w5, 
            w6=> c0_n49_w6, 
            w7=> c0_n49_w7, 
            w8=> c0_n49_w8, 
            w9=> c0_n49_w9, 
            w10=> c0_n49_w10, 
            w11=> c0_n49_w11, 
            w12=> c0_n49_w12, 
            w13=> c0_n49_w13, 
            w14=> c0_n49_w14, 
            w15=> c0_n49_w15, 
            w16=> c0_n49_w16, 
            w17=> c0_n49_w17, 
            w18=> c0_n49_w18, 
            w19=> c0_n49_w19, 
            w20=> c0_n49_w20, 
            w21=> c0_n49_w21, 
            w22=> c0_n49_w22, 
            w23=> c0_n49_w23, 
            w24=> c0_n49_w24, 
            w25=> c0_n49_w25, 
            w26=> c0_n49_w26, 
            w27=> c0_n49_w27, 
            w28=> c0_n49_w28, 
            w29=> c0_n49_w29, 
            w30=> c0_n49_w30, 
            w31=> c0_n49_w31, 
            w32=> c0_n49_w32, 
            w33=> c0_n49_w33, 
            w34=> c0_n49_w34, 
            w35=> c0_n49_w35, 
            w36=> c0_n49_w36, 
            w37=> c0_n49_w37, 
            w38=> c0_n49_w38, 
            w39=> c0_n49_w39, 
            w40=> c0_n49_w40, 
            w41=> c0_n49_w41, 
            w42=> c0_n49_w42, 
            w43=> c0_n49_w43, 
            w44=> c0_n49_w44, 
            w45=> c0_n49_w45, 
            w46=> c0_n49_w46, 
            w47=> c0_n49_w47, 
            w48=> c0_n49_w48, 
            w49=> c0_n49_w49, 
            w50=> c0_n49_w50, 
            w51=> c0_n49_w51, 
            w52=> c0_n49_w52, 
            w53=> c0_n49_w53, 
            w54=> c0_n49_w54, 
            w55=> c0_n49_w55, 
            w56=> c0_n49_w56, 
            w57=> c0_n49_w57, 
            w58=> c0_n49_w58, 
            w59=> c0_n49_w59, 
            w60=> c0_n49_w60, 
            w61=> c0_n49_w61, 
            w62=> c0_n49_w62, 
            w63=> c0_n49_w63, 
            w64=> c0_n49_w64, 
            w65=> c0_n49_w65, 
            w66=> c0_n49_w66, 
            w67=> c0_n49_w67, 
            w68=> c0_n49_w68, 
            w69=> c0_n49_w69, 
            w70=> c0_n49_w70, 
            w71=> c0_n49_w71, 
            w72=> c0_n49_w72, 
            w73=> c0_n49_w73, 
            w74=> c0_n49_w74, 
            w75=> c0_n49_w75, 
            w76=> c0_n49_w76, 
            w77=> c0_n49_w77, 
            w78=> c0_n49_w78, 
            w79=> c0_n49_w79, 
            w80=> c0_n49_w80, 
            w81=> c0_n49_w81, 
            w82=> c0_n49_w82, 
            w83=> c0_n49_w83, 
            w84=> c0_n49_w84, 
            w85=> c0_n49_w85, 
            w86=> c0_n49_w86, 
            w87=> c0_n49_w87, 
            w88=> c0_n49_w88, 
            w89=> c0_n49_w89, 
            w90=> c0_n49_w90, 
            w91=> c0_n49_w91, 
            w92=> c0_n49_w92, 
            w93=> c0_n49_w93, 
            w94=> c0_n49_w94, 
            w95=> c0_n49_w95, 
            w96=> c0_n49_w96, 
            w97=> c0_n49_w97, 
            w98=> c0_n49_w98, 
            w99=> c0_n49_w99, 
            w100=> c0_n49_w100, 
            w101=> c0_n49_w101, 
            w102=> c0_n49_w102, 
            w103=> c0_n49_w103, 
            w104=> c0_n49_w104, 
            w105=> c0_n49_w105, 
            w106=> c0_n49_w106, 
            w107=> c0_n49_w107, 
            w108=> c0_n49_w108, 
            w109=> c0_n49_w109, 
            w110=> c0_n49_w110, 
            w111=> c0_n49_w111, 
            w112=> c0_n49_w112, 
            w113=> c0_n49_w113, 
            w114=> c0_n49_w114, 
            w115=> c0_n49_w115, 
            w116=> c0_n49_w116, 
            w117=> c0_n49_w117, 
            w118=> c0_n49_w118, 
            w119=> c0_n49_w119, 
            w120=> c0_n49_w120, 
            w121=> c0_n49_w121, 
            w122=> c0_n49_w122, 
            w123=> c0_n49_w123, 
            w124=> c0_n49_w124, 
            w125=> c0_n49_w125, 
            w126=> c0_n49_w126, 
            w127=> c0_n49_w127, 
            w128=> c0_n49_w128, 
            w129=> c0_n49_w129, 
            w130=> c0_n49_w130, 
            w131=> c0_n49_w131, 
            w132=> c0_n49_w132, 
            w133=> c0_n49_w133, 
            w134=> c0_n49_w134, 
            w135=> c0_n49_w135, 
            w136=> c0_n49_w136, 
            w137=> c0_n49_w137, 
            w138=> c0_n49_w138, 
            w139=> c0_n49_w139, 
            w140=> c0_n49_w140, 
            w141=> c0_n49_w141, 
            w142=> c0_n49_w142, 
            w143=> c0_n49_w143, 
            w144=> c0_n49_w144, 
            w145=> c0_n49_w145, 
            w146=> c0_n49_w146, 
            w147=> c0_n49_w147, 
            w148=> c0_n49_w148, 
            w149=> c0_n49_w149, 
            w150=> c0_n49_w150, 
            w151=> c0_n49_w151, 
            w152=> c0_n49_w152, 
            w153=> c0_n49_w153, 
            w154=> c0_n49_w154, 
            w155=> c0_n49_w155, 
            w156=> c0_n49_w156, 
            w157=> c0_n49_w157, 
            w158=> c0_n49_w158, 
            w159=> c0_n49_w159, 
            w160=> c0_n49_w160, 
            w161=> c0_n49_w161, 
            w162=> c0_n49_w162, 
            w163=> c0_n49_w163, 
            w164=> c0_n49_w164, 
            w165=> c0_n49_w165, 
            w166=> c0_n49_w166, 
            w167=> c0_n49_w167, 
            w168=> c0_n49_w168, 
            w169=> c0_n49_w169, 
            w170=> c0_n49_w170, 
            w171=> c0_n49_w171, 
            w172=> c0_n49_w172, 
            w173=> c0_n49_w173, 
            w174=> c0_n49_w174, 
            w175=> c0_n49_w175, 
            w176=> c0_n49_w176, 
            w177=> c0_n49_w177, 
            w178=> c0_n49_w178, 
            w179=> c0_n49_w179, 
            w180=> c0_n49_w180, 
            w181=> c0_n49_w181, 
            w182=> c0_n49_w182, 
            w183=> c0_n49_w183, 
            w184=> c0_n49_w184, 
            w185=> c0_n49_w185, 
            w186=> c0_n49_w186, 
            w187=> c0_n49_w187, 
            w188=> c0_n49_w188, 
            w189=> c0_n49_w189, 
            w190=> c0_n49_w190, 
            w191=> c0_n49_w191, 
            w192=> c0_n49_w192, 
            w193=> c0_n49_w193, 
            w194=> c0_n49_w194, 
            w195=> c0_n49_w195, 
            w196=> c0_n49_w196, 
            w197=> c0_n49_w197, 
            w198=> c0_n49_w198, 
            w199=> c0_n49_w199, 
            w200=> c0_n49_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n49_y
   );           
            
neuron_inst_50: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n50_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n50_w1, 
            w2=> c0_n50_w2, 
            w3=> c0_n50_w3, 
            w4=> c0_n50_w4, 
            w5=> c0_n50_w5, 
            w6=> c0_n50_w6, 
            w7=> c0_n50_w7, 
            w8=> c0_n50_w8, 
            w9=> c0_n50_w9, 
            w10=> c0_n50_w10, 
            w11=> c0_n50_w11, 
            w12=> c0_n50_w12, 
            w13=> c0_n50_w13, 
            w14=> c0_n50_w14, 
            w15=> c0_n50_w15, 
            w16=> c0_n50_w16, 
            w17=> c0_n50_w17, 
            w18=> c0_n50_w18, 
            w19=> c0_n50_w19, 
            w20=> c0_n50_w20, 
            w21=> c0_n50_w21, 
            w22=> c0_n50_w22, 
            w23=> c0_n50_w23, 
            w24=> c0_n50_w24, 
            w25=> c0_n50_w25, 
            w26=> c0_n50_w26, 
            w27=> c0_n50_w27, 
            w28=> c0_n50_w28, 
            w29=> c0_n50_w29, 
            w30=> c0_n50_w30, 
            w31=> c0_n50_w31, 
            w32=> c0_n50_w32, 
            w33=> c0_n50_w33, 
            w34=> c0_n50_w34, 
            w35=> c0_n50_w35, 
            w36=> c0_n50_w36, 
            w37=> c0_n50_w37, 
            w38=> c0_n50_w38, 
            w39=> c0_n50_w39, 
            w40=> c0_n50_w40, 
            w41=> c0_n50_w41, 
            w42=> c0_n50_w42, 
            w43=> c0_n50_w43, 
            w44=> c0_n50_w44, 
            w45=> c0_n50_w45, 
            w46=> c0_n50_w46, 
            w47=> c0_n50_w47, 
            w48=> c0_n50_w48, 
            w49=> c0_n50_w49, 
            w50=> c0_n50_w50, 
            w51=> c0_n50_w51, 
            w52=> c0_n50_w52, 
            w53=> c0_n50_w53, 
            w54=> c0_n50_w54, 
            w55=> c0_n50_w55, 
            w56=> c0_n50_w56, 
            w57=> c0_n50_w57, 
            w58=> c0_n50_w58, 
            w59=> c0_n50_w59, 
            w60=> c0_n50_w60, 
            w61=> c0_n50_w61, 
            w62=> c0_n50_w62, 
            w63=> c0_n50_w63, 
            w64=> c0_n50_w64, 
            w65=> c0_n50_w65, 
            w66=> c0_n50_w66, 
            w67=> c0_n50_w67, 
            w68=> c0_n50_w68, 
            w69=> c0_n50_w69, 
            w70=> c0_n50_w70, 
            w71=> c0_n50_w71, 
            w72=> c0_n50_w72, 
            w73=> c0_n50_w73, 
            w74=> c0_n50_w74, 
            w75=> c0_n50_w75, 
            w76=> c0_n50_w76, 
            w77=> c0_n50_w77, 
            w78=> c0_n50_w78, 
            w79=> c0_n50_w79, 
            w80=> c0_n50_w80, 
            w81=> c0_n50_w81, 
            w82=> c0_n50_w82, 
            w83=> c0_n50_w83, 
            w84=> c0_n50_w84, 
            w85=> c0_n50_w85, 
            w86=> c0_n50_w86, 
            w87=> c0_n50_w87, 
            w88=> c0_n50_w88, 
            w89=> c0_n50_w89, 
            w90=> c0_n50_w90, 
            w91=> c0_n50_w91, 
            w92=> c0_n50_w92, 
            w93=> c0_n50_w93, 
            w94=> c0_n50_w94, 
            w95=> c0_n50_w95, 
            w96=> c0_n50_w96, 
            w97=> c0_n50_w97, 
            w98=> c0_n50_w98, 
            w99=> c0_n50_w99, 
            w100=> c0_n50_w100, 
            w101=> c0_n50_w101, 
            w102=> c0_n50_w102, 
            w103=> c0_n50_w103, 
            w104=> c0_n50_w104, 
            w105=> c0_n50_w105, 
            w106=> c0_n50_w106, 
            w107=> c0_n50_w107, 
            w108=> c0_n50_w108, 
            w109=> c0_n50_w109, 
            w110=> c0_n50_w110, 
            w111=> c0_n50_w111, 
            w112=> c0_n50_w112, 
            w113=> c0_n50_w113, 
            w114=> c0_n50_w114, 
            w115=> c0_n50_w115, 
            w116=> c0_n50_w116, 
            w117=> c0_n50_w117, 
            w118=> c0_n50_w118, 
            w119=> c0_n50_w119, 
            w120=> c0_n50_w120, 
            w121=> c0_n50_w121, 
            w122=> c0_n50_w122, 
            w123=> c0_n50_w123, 
            w124=> c0_n50_w124, 
            w125=> c0_n50_w125, 
            w126=> c0_n50_w126, 
            w127=> c0_n50_w127, 
            w128=> c0_n50_w128, 
            w129=> c0_n50_w129, 
            w130=> c0_n50_w130, 
            w131=> c0_n50_w131, 
            w132=> c0_n50_w132, 
            w133=> c0_n50_w133, 
            w134=> c0_n50_w134, 
            w135=> c0_n50_w135, 
            w136=> c0_n50_w136, 
            w137=> c0_n50_w137, 
            w138=> c0_n50_w138, 
            w139=> c0_n50_w139, 
            w140=> c0_n50_w140, 
            w141=> c0_n50_w141, 
            w142=> c0_n50_w142, 
            w143=> c0_n50_w143, 
            w144=> c0_n50_w144, 
            w145=> c0_n50_w145, 
            w146=> c0_n50_w146, 
            w147=> c0_n50_w147, 
            w148=> c0_n50_w148, 
            w149=> c0_n50_w149, 
            w150=> c0_n50_w150, 
            w151=> c0_n50_w151, 
            w152=> c0_n50_w152, 
            w153=> c0_n50_w153, 
            w154=> c0_n50_w154, 
            w155=> c0_n50_w155, 
            w156=> c0_n50_w156, 
            w157=> c0_n50_w157, 
            w158=> c0_n50_w158, 
            w159=> c0_n50_w159, 
            w160=> c0_n50_w160, 
            w161=> c0_n50_w161, 
            w162=> c0_n50_w162, 
            w163=> c0_n50_w163, 
            w164=> c0_n50_w164, 
            w165=> c0_n50_w165, 
            w166=> c0_n50_w166, 
            w167=> c0_n50_w167, 
            w168=> c0_n50_w168, 
            w169=> c0_n50_w169, 
            w170=> c0_n50_w170, 
            w171=> c0_n50_w171, 
            w172=> c0_n50_w172, 
            w173=> c0_n50_w173, 
            w174=> c0_n50_w174, 
            w175=> c0_n50_w175, 
            w176=> c0_n50_w176, 
            w177=> c0_n50_w177, 
            w178=> c0_n50_w178, 
            w179=> c0_n50_w179, 
            w180=> c0_n50_w180, 
            w181=> c0_n50_w181, 
            w182=> c0_n50_w182, 
            w183=> c0_n50_w183, 
            w184=> c0_n50_w184, 
            w185=> c0_n50_w185, 
            w186=> c0_n50_w186, 
            w187=> c0_n50_w187, 
            w188=> c0_n50_w188, 
            w189=> c0_n50_w189, 
            w190=> c0_n50_w190, 
            w191=> c0_n50_w191, 
            w192=> c0_n50_w192, 
            w193=> c0_n50_w193, 
            w194=> c0_n50_w194, 
            w195=> c0_n50_w195, 
            w196=> c0_n50_w196, 
            w197=> c0_n50_w197, 
            w198=> c0_n50_w198, 
            w199=> c0_n50_w199, 
            w200=> c0_n50_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n50_y
   );           
            
neuron_inst_51: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n51_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n51_w1, 
            w2=> c0_n51_w2, 
            w3=> c0_n51_w3, 
            w4=> c0_n51_w4, 
            w5=> c0_n51_w5, 
            w6=> c0_n51_w6, 
            w7=> c0_n51_w7, 
            w8=> c0_n51_w8, 
            w9=> c0_n51_w9, 
            w10=> c0_n51_w10, 
            w11=> c0_n51_w11, 
            w12=> c0_n51_w12, 
            w13=> c0_n51_w13, 
            w14=> c0_n51_w14, 
            w15=> c0_n51_w15, 
            w16=> c0_n51_w16, 
            w17=> c0_n51_w17, 
            w18=> c0_n51_w18, 
            w19=> c0_n51_w19, 
            w20=> c0_n51_w20, 
            w21=> c0_n51_w21, 
            w22=> c0_n51_w22, 
            w23=> c0_n51_w23, 
            w24=> c0_n51_w24, 
            w25=> c0_n51_w25, 
            w26=> c0_n51_w26, 
            w27=> c0_n51_w27, 
            w28=> c0_n51_w28, 
            w29=> c0_n51_w29, 
            w30=> c0_n51_w30, 
            w31=> c0_n51_w31, 
            w32=> c0_n51_w32, 
            w33=> c0_n51_w33, 
            w34=> c0_n51_w34, 
            w35=> c0_n51_w35, 
            w36=> c0_n51_w36, 
            w37=> c0_n51_w37, 
            w38=> c0_n51_w38, 
            w39=> c0_n51_w39, 
            w40=> c0_n51_w40, 
            w41=> c0_n51_w41, 
            w42=> c0_n51_w42, 
            w43=> c0_n51_w43, 
            w44=> c0_n51_w44, 
            w45=> c0_n51_w45, 
            w46=> c0_n51_w46, 
            w47=> c0_n51_w47, 
            w48=> c0_n51_w48, 
            w49=> c0_n51_w49, 
            w50=> c0_n51_w50, 
            w51=> c0_n51_w51, 
            w52=> c0_n51_w52, 
            w53=> c0_n51_w53, 
            w54=> c0_n51_w54, 
            w55=> c0_n51_w55, 
            w56=> c0_n51_w56, 
            w57=> c0_n51_w57, 
            w58=> c0_n51_w58, 
            w59=> c0_n51_w59, 
            w60=> c0_n51_w60, 
            w61=> c0_n51_w61, 
            w62=> c0_n51_w62, 
            w63=> c0_n51_w63, 
            w64=> c0_n51_w64, 
            w65=> c0_n51_w65, 
            w66=> c0_n51_w66, 
            w67=> c0_n51_w67, 
            w68=> c0_n51_w68, 
            w69=> c0_n51_w69, 
            w70=> c0_n51_w70, 
            w71=> c0_n51_w71, 
            w72=> c0_n51_w72, 
            w73=> c0_n51_w73, 
            w74=> c0_n51_w74, 
            w75=> c0_n51_w75, 
            w76=> c0_n51_w76, 
            w77=> c0_n51_w77, 
            w78=> c0_n51_w78, 
            w79=> c0_n51_w79, 
            w80=> c0_n51_w80, 
            w81=> c0_n51_w81, 
            w82=> c0_n51_w82, 
            w83=> c0_n51_w83, 
            w84=> c0_n51_w84, 
            w85=> c0_n51_w85, 
            w86=> c0_n51_w86, 
            w87=> c0_n51_w87, 
            w88=> c0_n51_w88, 
            w89=> c0_n51_w89, 
            w90=> c0_n51_w90, 
            w91=> c0_n51_w91, 
            w92=> c0_n51_w92, 
            w93=> c0_n51_w93, 
            w94=> c0_n51_w94, 
            w95=> c0_n51_w95, 
            w96=> c0_n51_w96, 
            w97=> c0_n51_w97, 
            w98=> c0_n51_w98, 
            w99=> c0_n51_w99, 
            w100=> c0_n51_w100, 
            w101=> c0_n51_w101, 
            w102=> c0_n51_w102, 
            w103=> c0_n51_w103, 
            w104=> c0_n51_w104, 
            w105=> c0_n51_w105, 
            w106=> c0_n51_w106, 
            w107=> c0_n51_w107, 
            w108=> c0_n51_w108, 
            w109=> c0_n51_w109, 
            w110=> c0_n51_w110, 
            w111=> c0_n51_w111, 
            w112=> c0_n51_w112, 
            w113=> c0_n51_w113, 
            w114=> c0_n51_w114, 
            w115=> c0_n51_w115, 
            w116=> c0_n51_w116, 
            w117=> c0_n51_w117, 
            w118=> c0_n51_w118, 
            w119=> c0_n51_w119, 
            w120=> c0_n51_w120, 
            w121=> c0_n51_w121, 
            w122=> c0_n51_w122, 
            w123=> c0_n51_w123, 
            w124=> c0_n51_w124, 
            w125=> c0_n51_w125, 
            w126=> c0_n51_w126, 
            w127=> c0_n51_w127, 
            w128=> c0_n51_w128, 
            w129=> c0_n51_w129, 
            w130=> c0_n51_w130, 
            w131=> c0_n51_w131, 
            w132=> c0_n51_w132, 
            w133=> c0_n51_w133, 
            w134=> c0_n51_w134, 
            w135=> c0_n51_w135, 
            w136=> c0_n51_w136, 
            w137=> c0_n51_w137, 
            w138=> c0_n51_w138, 
            w139=> c0_n51_w139, 
            w140=> c0_n51_w140, 
            w141=> c0_n51_w141, 
            w142=> c0_n51_w142, 
            w143=> c0_n51_w143, 
            w144=> c0_n51_w144, 
            w145=> c0_n51_w145, 
            w146=> c0_n51_w146, 
            w147=> c0_n51_w147, 
            w148=> c0_n51_w148, 
            w149=> c0_n51_w149, 
            w150=> c0_n51_w150, 
            w151=> c0_n51_w151, 
            w152=> c0_n51_w152, 
            w153=> c0_n51_w153, 
            w154=> c0_n51_w154, 
            w155=> c0_n51_w155, 
            w156=> c0_n51_w156, 
            w157=> c0_n51_w157, 
            w158=> c0_n51_w158, 
            w159=> c0_n51_w159, 
            w160=> c0_n51_w160, 
            w161=> c0_n51_w161, 
            w162=> c0_n51_w162, 
            w163=> c0_n51_w163, 
            w164=> c0_n51_w164, 
            w165=> c0_n51_w165, 
            w166=> c0_n51_w166, 
            w167=> c0_n51_w167, 
            w168=> c0_n51_w168, 
            w169=> c0_n51_w169, 
            w170=> c0_n51_w170, 
            w171=> c0_n51_w171, 
            w172=> c0_n51_w172, 
            w173=> c0_n51_w173, 
            w174=> c0_n51_w174, 
            w175=> c0_n51_w175, 
            w176=> c0_n51_w176, 
            w177=> c0_n51_w177, 
            w178=> c0_n51_w178, 
            w179=> c0_n51_w179, 
            w180=> c0_n51_w180, 
            w181=> c0_n51_w181, 
            w182=> c0_n51_w182, 
            w183=> c0_n51_w183, 
            w184=> c0_n51_w184, 
            w185=> c0_n51_w185, 
            w186=> c0_n51_w186, 
            w187=> c0_n51_w187, 
            w188=> c0_n51_w188, 
            w189=> c0_n51_w189, 
            w190=> c0_n51_w190, 
            w191=> c0_n51_w191, 
            w192=> c0_n51_w192, 
            w193=> c0_n51_w193, 
            w194=> c0_n51_w194, 
            w195=> c0_n51_w195, 
            w196=> c0_n51_w196, 
            w197=> c0_n51_w197, 
            w198=> c0_n51_w198, 
            w199=> c0_n51_w199, 
            w200=> c0_n51_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n51_y
   );           
            
neuron_inst_52: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n52_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n52_w1, 
            w2=> c0_n52_w2, 
            w3=> c0_n52_w3, 
            w4=> c0_n52_w4, 
            w5=> c0_n52_w5, 
            w6=> c0_n52_w6, 
            w7=> c0_n52_w7, 
            w8=> c0_n52_w8, 
            w9=> c0_n52_w9, 
            w10=> c0_n52_w10, 
            w11=> c0_n52_w11, 
            w12=> c0_n52_w12, 
            w13=> c0_n52_w13, 
            w14=> c0_n52_w14, 
            w15=> c0_n52_w15, 
            w16=> c0_n52_w16, 
            w17=> c0_n52_w17, 
            w18=> c0_n52_w18, 
            w19=> c0_n52_w19, 
            w20=> c0_n52_w20, 
            w21=> c0_n52_w21, 
            w22=> c0_n52_w22, 
            w23=> c0_n52_w23, 
            w24=> c0_n52_w24, 
            w25=> c0_n52_w25, 
            w26=> c0_n52_w26, 
            w27=> c0_n52_w27, 
            w28=> c0_n52_w28, 
            w29=> c0_n52_w29, 
            w30=> c0_n52_w30, 
            w31=> c0_n52_w31, 
            w32=> c0_n52_w32, 
            w33=> c0_n52_w33, 
            w34=> c0_n52_w34, 
            w35=> c0_n52_w35, 
            w36=> c0_n52_w36, 
            w37=> c0_n52_w37, 
            w38=> c0_n52_w38, 
            w39=> c0_n52_w39, 
            w40=> c0_n52_w40, 
            w41=> c0_n52_w41, 
            w42=> c0_n52_w42, 
            w43=> c0_n52_w43, 
            w44=> c0_n52_w44, 
            w45=> c0_n52_w45, 
            w46=> c0_n52_w46, 
            w47=> c0_n52_w47, 
            w48=> c0_n52_w48, 
            w49=> c0_n52_w49, 
            w50=> c0_n52_w50, 
            w51=> c0_n52_w51, 
            w52=> c0_n52_w52, 
            w53=> c0_n52_w53, 
            w54=> c0_n52_w54, 
            w55=> c0_n52_w55, 
            w56=> c0_n52_w56, 
            w57=> c0_n52_w57, 
            w58=> c0_n52_w58, 
            w59=> c0_n52_w59, 
            w60=> c0_n52_w60, 
            w61=> c0_n52_w61, 
            w62=> c0_n52_w62, 
            w63=> c0_n52_w63, 
            w64=> c0_n52_w64, 
            w65=> c0_n52_w65, 
            w66=> c0_n52_w66, 
            w67=> c0_n52_w67, 
            w68=> c0_n52_w68, 
            w69=> c0_n52_w69, 
            w70=> c0_n52_w70, 
            w71=> c0_n52_w71, 
            w72=> c0_n52_w72, 
            w73=> c0_n52_w73, 
            w74=> c0_n52_w74, 
            w75=> c0_n52_w75, 
            w76=> c0_n52_w76, 
            w77=> c0_n52_w77, 
            w78=> c0_n52_w78, 
            w79=> c0_n52_w79, 
            w80=> c0_n52_w80, 
            w81=> c0_n52_w81, 
            w82=> c0_n52_w82, 
            w83=> c0_n52_w83, 
            w84=> c0_n52_w84, 
            w85=> c0_n52_w85, 
            w86=> c0_n52_w86, 
            w87=> c0_n52_w87, 
            w88=> c0_n52_w88, 
            w89=> c0_n52_w89, 
            w90=> c0_n52_w90, 
            w91=> c0_n52_w91, 
            w92=> c0_n52_w92, 
            w93=> c0_n52_w93, 
            w94=> c0_n52_w94, 
            w95=> c0_n52_w95, 
            w96=> c0_n52_w96, 
            w97=> c0_n52_w97, 
            w98=> c0_n52_w98, 
            w99=> c0_n52_w99, 
            w100=> c0_n52_w100, 
            w101=> c0_n52_w101, 
            w102=> c0_n52_w102, 
            w103=> c0_n52_w103, 
            w104=> c0_n52_w104, 
            w105=> c0_n52_w105, 
            w106=> c0_n52_w106, 
            w107=> c0_n52_w107, 
            w108=> c0_n52_w108, 
            w109=> c0_n52_w109, 
            w110=> c0_n52_w110, 
            w111=> c0_n52_w111, 
            w112=> c0_n52_w112, 
            w113=> c0_n52_w113, 
            w114=> c0_n52_w114, 
            w115=> c0_n52_w115, 
            w116=> c0_n52_w116, 
            w117=> c0_n52_w117, 
            w118=> c0_n52_w118, 
            w119=> c0_n52_w119, 
            w120=> c0_n52_w120, 
            w121=> c0_n52_w121, 
            w122=> c0_n52_w122, 
            w123=> c0_n52_w123, 
            w124=> c0_n52_w124, 
            w125=> c0_n52_w125, 
            w126=> c0_n52_w126, 
            w127=> c0_n52_w127, 
            w128=> c0_n52_w128, 
            w129=> c0_n52_w129, 
            w130=> c0_n52_w130, 
            w131=> c0_n52_w131, 
            w132=> c0_n52_w132, 
            w133=> c0_n52_w133, 
            w134=> c0_n52_w134, 
            w135=> c0_n52_w135, 
            w136=> c0_n52_w136, 
            w137=> c0_n52_w137, 
            w138=> c0_n52_w138, 
            w139=> c0_n52_w139, 
            w140=> c0_n52_w140, 
            w141=> c0_n52_w141, 
            w142=> c0_n52_w142, 
            w143=> c0_n52_w143, 
            w144=> c0_n52_w144, 
            w145=> c0_n52_w145, 
            w146=> c0_n52_w146, 
            w147=> c0_n52_w147, 
            w148=> c0_n52_w148, 
            w149=> c0_n52_w149, 
            w150=> c0_n52_w150, 
            w151=> c0_n52_w151, 
            w152=> c0_n52_w152, 
            w153=> c0_n52_w153, 
            w154=> c0_n52_w154, 
            w155=> c0_n52_w155, 
            w156=> c0_n52_w156, 
            w157=> c0_n52_w157, 
            w158=> c0_n52_w158, 
            w159=> c0_n52_w159, 
            w160=> c0_n52_w160, 
            w161=> c0_n52_w161, 
            w162=> c0_n52_w162, 
            w163=> c0_n52_w163, 
            w164=> c0_n52_w164, 
            w165=> c0_n52_w165, 
            w166=> c0_n52_w166, 
            w167=> c0_n52_w167, 
            w168=> c0_n52_w168, 
            w169=> c0_n52_w169, 
            w170=> c0_n52_w170, 
            w171=> c0_n52_w171, 
            w172=> c0_n52_w172, 
            w173=> c0_n52_w173, 
            w174=> c0_n52_w174, 
            w175=> c0_n52_w175, 
            w176=> c0_n52_w176, 
            w177=> c0_n52_w177, 
            w178=> c0_n52_w178, 
            w179=> c0_n52_w179, 
            w180=> c0_n52_w180, 
            w181=> c0_n52_w181, 
            w182=> c0_n52_w182, 
            w183=> c0_n52_w183, 
            w184=> c0_n52_w184, 
            w185=> c0_n52_w185, 
            w186=> c0_n52_w186, 
            w187=> c0_n52_w187, 
            w188=> c0_n52_w188, 
            w189=> c0_n52_w189, 
            w190=> c0_n52_w190, 
            w191=> c0_n52_w191, 
            w192=> c0_n52_w192, 
            w193=> c0_n52_w193, 
            w194=> c0_n52_w194, 
            w195=> c0_n52_w195, 
            w196=> c0_n52_w196, 
            w197=> c0_n52_w197, 
            w198=> c0_n52_w198, 
            w199=> c0_n52_w199, 
            w200=> c0_n52_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n52_y
   );           
            
neuron_inst_53: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n53_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n53_w1, 
            w2=> c0_n53_w2, 
            w3=> c0_n53_w3, 
            w4=> c0_n53_w4, 
            w5=> c0_n53_w5, 
            w6=> c0_n53_w6, 
            w7=> c0_n53_w7, 
            w8=> c0_n53_w8, 
            w9=> c0_n53_w9, 
            w10=> c0_n53_w10, 
            w11=> c0_n53_w11, 
            w12=> c0_n53_w12, 
            w13=> c0_n53_w13, 
            w14=> c0_n53_w14, 
            w15=> c0_n53_w15, 
            w16=> c0_n53_w16, 
            w17=> c0_n53_w17, 
            w18=> c0_n53_w18, 
            w19=> c0_n53_w19, 
            w20=> c0_n53_w20, 
            w21=> c0_n53_w21, 
            w22=> c0_n53_w22, 
            w23=> c0_n53_w23, 
            w24=> c0_n53_w24, 
            w25=> c0_n53_w25, 
            w26=> c0_n53_w26, 
            w27=> c0_n53_w27, 
            w28=> c0_n53_w28, 
            w29=> c0_n53_w29, 
            w30=> c0_n53_w30, 
            w31=> c0_n53_w31, 
            w32=> c0_n53_w32, 
            w33=> c0_n53_w33, 
            w34=> c0_n53_w34, 
            w35=> c0_n53_w35, 
            w36=> c0_n53_w36, 
            w37=> c0_n53_w37, 
            w38=> c0_n53_w38, 
            w39=> c0_n53_w39, 
            w40=> c0_n53_w40, 
            w41=> c0_n53_w41, 
            w42=> c0_n53_w42, 
            w43=> c0_n53_w43, 
            w44=> c0_n53_w44, 
            w45=> c0_n53_w45, 
            w46=> c0_n53_w46, 
            w47=> c0_n53_w47, 
            w48=> c0_n53_w48, 
            w49=> c0_n53_w49, 
            w50=> c0_n53_w50, 
            w51=> c0_n53_w51, 
            w52=> c0_n53_w52, 
            w53=> c0_n53_w53, 
            w54=> c0_n53_w54, 
            w55=> c0_n53_w55, 
            w56=> c0_n53_w56, 
            w57=> c0_n53_w57, 
            w58=> c0_n53_w58, 
            w59=> c0_n53_w59, 
            w60=> c0_n53_w60, 
            w61=> c0_n53_w61, 
            w62=> c0_n53_w62, 
            w63=> c0_n53_w63, 
            w64=> c0_n53_w64, 
            w65=> c0_n53_w65, 
            w66=> c0_n53_w66, 
            w67=> c0_n53_w67, 
            w68=> c0_n53_w68, 
            w69=> c0_n53_w69, 
            w70=> c0_n53_w70, 
            w71=> c0_n53_w71, 
            w72=> c0_n53_w72, 
            w73=> c0_n53_w73, 
            w74=> c0_n53_w74, 
            w75=> c0_n53_w75, 
            w76=> c0_n53_w76, 
            w77=> c0_n53_w77, 
            w78=> c0_n53_w78, 
            w79=> c0_n53_w79, 
            w80=> c0_n53_w80, 
            w81=> c0_n53_w81, 
            w82=> c0_n53_w82, 
            w83=> c0_n53_w83, 
            w84=> c0_n53_w84, 
            w85=> c0_n53_w85, 
            w86=> c0_n53_w86, 
            w87=> c0_n53_w87, 
            w88=> c0_n53_w88, 
            w89=> c0_n53_w89, 
            w90=> c0_n53_w90, 
            w91=> c0_n53_w91, 
            w92=> c0_n53_w92, 
            w93=> c0_n53_w93, 
            w94=> c0_n53_w94, 
            w95=> c0_n53_w95, 
            w96=> c0_n53_w96, 
            w97=> c0_n53_w97, 
            w98=> c0_n53_w98, 
            w99=> c0_n53_w99, 
            w100=> c0_n53_w100, 
            w101=> c0_n53_w101, 
            w102=> c0_n53_w102, 
            w103=> c0_n53_w103, 
            w104=> c0_n53_w104, 
            w105=> c0_n53_w105, 
            w106=> c0_n53_w106, 
            w107=> c0_n53_w107, 
            w108=> c0_n53_w108, 
            w109=> c0_n53_w109, 
            w110=> c0_n53_w110, 
            w111=> c0_n53_w111, 
            w112=> c0_n53_w112, 
            w113=> c0_n53_w113, 
            w114=> c0_n53_w114, 
            w115=> c0_n53_w115, 
            w116=> c0_n53_w116, 
            w117=> c0_n53_w117, 
            w118=> c0_n53_w118, 
            w119=> c0_n53_w119, 
            w120=> c0_n53_w120, 
            w121=> c0_n53_w121, 
            w122=> c0_n53_w122, 
            w123=> c0_n53_w123, 
            w124=> c0_n53_w124, 
            w125=> c0_n53_w125, 
            w126=> c0_n53_w126, 
            w127=> c0_n53_w127, 
            w128=> c0_n53_w128, 
            w129=> c0_n53_w129, 
            w130=> c0_n53_w130, 
            w131=> c0_n53_w131, 
            w132=> c0_n53_w132, 
            w133=> c0_n53_w133, 
            w134=> c0_n53_w134, 
            w135=> c0_n53_w135, 
            w136=> c0_n53_w136, 
            w137=> c0_n53_w137, 
            w138=> c0_n53_w138, 
            w139=> c0_n53_w139, 
            w140=> c0_n53_w140, 
            w141=> c0_n53_w141, 
            w142=> c0_n53_w142, 
            w143=> c0_n53_w143, 
            w144=> c0_n53_w144, 
            w145=> c0_n53_w145, 
            w146=> c0_n53_w146, 
            w147=> c0_n53_w147, 
            w148=> c0_n53_w148, 
            w149=> c0_n53_w149, 
            w150=> c0_n53_w150, 
            w151=> c0_n53_w151, 
            w152=> c0_n53_w152, 
            w153=> c0_n53_w153, 
            w154=> c0_n53_w154, 
            w155=> c0_n53_w155, 
            w156=> c0_n53_w156, 
            w157=> c0_n53_w157, 
            w158=> c0_n53_w158, 
            w159=> c0_n53_w159, 
            w160=> c0_n53_w160, 
            w161=> c0_n53_w161, 
            w162=> c0_n53_w162, 
            w163=> c0_n53_w163, 
            w164=> c0_n53_w164, 
            w165=> c0_n53_w165, 
            w166=> c0_n53_w166, 
            w167=> c0_n53_w167, 
            w168=> c0_n53_w168, 
            w169=> c0_n53_w169, 
            w170=> c0_n53_w170, 
            w171=> c0_n53_w171, 
            w172=> c0_n53_w172, 
            w173=> c0_n53_w173, 
            w174=> c0_n53_w174, 
            w175=> c0_n53_w175, 
            w176=> c0_n53_w176, 
            w177=> c0_n53_w177, 
            w178=> c0_n53_w178, 
            w179=> c0_n53_w179, 
            w180=> c0_n53_w180, 
            w181=> c0_n53_w181, 
            w182=> c0_n53_w182, 
            w183=> c0_n53_w183, 
            w184=> c0_n53_w184, 
            w185=> c0_n53_w185, 
            w186=> c0_n53_w186, 
            w187=> c0_n53_w187, 
            w188=> c0_n53_w188, 
            w189=> c0_n53_w189, 
            w190=> c0_n53_w190, 
            w191=> c0_n53_w191, 
            w192=> c0_n53_w192, 
            w193=> c0_n53_w193, 
            w194=> c0_n53_w194, 
            w195=> c0_n53_w195, 
            w196=> c0_n53_w196, 
            w197=> c0_n53_w197, 
            w198=> c0_n53_w198, 
            w199=> c0_n53_w199, 
            w200=> c0_n53_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n53_y
   );           
            
neuron_inst_54: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n54_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n54_w1, 
            w2=> c0_n54_w2, 
            w3=> c0_n54_w3, 
            w4=> c0_n54_w4, 
            w5=> c0_n54_w5, 
            w6=> c0_n54_w6, 
            w7=> c0_n54_w7, 
            w8=> c0_n54_w8, 
            w9=> c0_n54_w9, 
            w10=> c0_n54_w10, 
            w11=> c0_n54_w11, 
            w12=> c0_n54_w12, 
            w13=> c0_n54_w13, 
            w14=> c0_n54_w14, 
            w15=> c0_n54_w15, 
            w16=> c0_n54_w16, 
            w17=> c0_n54_w17, 
            w18=> c0_n54_w18, 
            w19=> c0_n54_w19, 
            w20=> c0_n54_w20, 
            w21=> c0_n54_w21, 
            w22=> c0_n54_w22, 
            w23=> c0_n54_w23, 
            w24=> c0_n54_w24, 
            w25=> c0_n54_w25, 
            w26=> c0_n54_w26, 
            w27=> c0_n54_w27, 
            w28=> c0_n54_w28, 
            w29=> c0_n54_w29, 
            w30=> c0_n54_w30, 
            w31=> c0_n54_w31, 
            w32=> c0_n54_w32, 
            w33=> c0_n54_w33, 
            w34=> c0_n54_w34, 
            w35=> c0_n54_w35, 
            w36=> c0_n54_w36, 
            w37=> c0_n54_w37, 
            w38=> c0_n54_w38, 
            w39=> c0_n54_w39, 
            w40=> c0_n54_w40, 
            w41=> c0_n54_w41, 
            w42=> c0_n54_w42, 
            w43=> c0_n54_w43, 
            w44=> c0_n54_w44, 
            w45=> c0_n54_w45, 
            w46=> c0_n54_w46, 
            w47=> c0_n54_w47, 
            w48=> c0_n54_w48, 
            w49=> c0_n54_w49, 
            w50=> c0_n54_w50, 
            w51=> c0_n54_w51, 
            w52=> c0_n54_w52, 
            w53=> c0_n54_w53, 
            w54=> c0_n54_w54, 
            w55=> c0_n54_w55, 
            w56=> c0_n54_w56, 
            w57=> c0_n54_w57, 
            w58=> c0_n54_w58, 
            w59=> c0_n54_w59, 
            w60=> c0_n54_w60, 
            w61=> c0_n54_w61, 
            w62=> c0_n54_w62, 
            w63=> c0_n54_w63, 
            w64=> c0_n54_w64, 
            w65=> c0_n54_w65, 
            w66=> c0_n54_w66, 
            w67=> c0_n54_w67, 
            w68=> c0_n54_w68, 
            w69=> c0_n54_w69, 
            w70=> c0_n54_w70, 
            w71=> c0_n54_w71, 
            w72=> c0_n54_w72, 
            w73=> c0_n54_w73, 
            w74=> c0_n54_w74, 
            w75=> c0_n54_w75, 
            w76=> c0_n54_w76, 
            w77=> c0_n54_w77, 
            w78=> c0_n54_w78, 
            w79=> c0_n54_w79, 
            w80=> c0_n54_w80, 
            w81=> c0_n54_w81, 
            w82=> c0_n54_w82, 
            w83=> c0_n54_w83, 
            w84=> c0_n54_w84, 
            w85=> c0_n54_w85, 
            w86=> c0_n54_w86, 
            w87=> c0_n54_w87, 
            w88=> c0_n54_w88, 
            w89=> c0_n54_w89, 
            w90=> c0_n54_w90, 
            w91=> c0_n54_w91, 
            w92=> c0_n54_w92, 
            w93=> c0_n54_w93, 
            w94=> c0_n54_w94, 
            w95=> c0_n54_w95, 
            w96=> c0_n54_w96, 
            w97=> c0_n54_w97, 
            w98=> c0_n54_w98, 
            w99=> c0_n54_w99, 
            w100=> c0_n54_w100, 
            w101=> c0_n54_w101, 
            w102=> c0_n54_w102, 
            w103=> c0_n54_w103, 
            w104=> c0_n54_w104, 
            w105=> c0_n54_w105, 
            w106=> c0_n54_w106, 
            w107=> c0_n54_w107, 
            w108=> c0_n54_w108, 
            w109=> c0_n54_w109, 
            w110=> c0_n54_w110, 
            w111=> c0_n54_w111, 
            w112=> c0_n54_w112, 
            w113=> c0_n54_w113, 
            w114=> c0_n54_w114, 
            w115=> c0_n54_w115, 
            w116=> c0_n54_w116, 
            w117=> c0_n54_w117, 
            w118=> c0_n54_w118, 
            w119=> c0_n54_w119, 
            w120=> c0_n54_w120, 
            w121=> c0_n54_w121, 
            w122=> c0_n54_w122, 
            w123=> c0_n54_w123, 
            w124=> c0_n54_w124, 
            w125=> c0_n54_w125, 
            w126=> c0_n54_w126, 
            w127=> c0_n54_w127, 
            w128=> c0_n54_w128, 
            w129=> c0_n54_w129, 
            w130=> c0_n54_w130, 
            w131=> c0_n54_w131, 
            w132=> c0_n54_w132, 
            w133=> c0_n54_w133, 
            w134=> c0_n54_w134, 
            w135=> c0_n54_w135, 
            w136=> c0_n54_w136, 
            w137=> c0_n54_w137, 
            w138=> c0_n54_w138, 
            w139=> c0_n54_w139, 
            w140=> c0_n54_w140, 
            w141=> c0_n54_w141, 
            w142=> c0_n54_w142, 
            w143=> c0_n54_w143, 
            w144=> c0_n54_w144, 
            w145=> c0_n54_w145, 
            w146=> c0_n54_w146, 
            w147=> c0_n54_w147, 
            w148=> c0_n54_w148, 
            w149=> c0_n54_w149, 
            w150=> c0_n54_w150, 
            w151=> c0_n54_w151, 
            w152=> c0_n54_w152, 
            w153=> c0_n54_w153, 
            w154=> c0_n54_w154, 
            w155=> c0_n54_w155, 
            w156=> c0_n54_w156, 
            w157=> c0_n54_w157, 
            w158=> c0_n54_w158, 
            w159=> c0_n54_w159, 
            w160=> c0_n54_w160, 
            w161=> c0_n54_w161, 
            w162=> c0_n54_w162, 
            w163=> c0_n54_w163, 
            w164=> c0_n54_w164, 
            w165=> c0_n54_w165, 
            w166=> c0_n54_w166, 
            w167=> c0_n54_w167, 
            w168=> c0_n54_w168, 
            w169=> c0_n54_w169, 
            w170=> c0_n54_w170, 
            w171=> c0_n54_w171, 
            w172=> c0_n54_w172, 
            w173=> c0_n54_w173, 
            w174=> c0_n54_w174, 
            w175=> c0_n54_w175, 
            w176=> c0_n54_w176, 
            w177=> c0_n54_w177, 
            w178=> c0_n54_w178, 
            w179=> c0_n54_w179, 
            w180=> c0_n54_w180, 
            w181=> c0_n54_w181, 
            w182=> c0_n54_w182, 
            w183=> c0_n54_w183, 
            w184=> c0_n54_w184, 
            w185=> c0_n54_w185, 
            w186=> c0_n54_w186, 
            w187=> c0_n54_w187, 
            w188=> c0_n54_w188, 
            w189=> c0_n54_w189, 
            w190=> c0_n54_w190, 
            w191=> c0_n54_w191, 
            w192=> c0_n54_w192, 
            w193=> c0_n54_w193, 
            w194=> c0_n54_w194, 
            w195=> c0_n54_w195, 
            w196=> c0_n54_w196, 
            w197=> c0_n54_w197, 
            w198=> c0_n54_w198, 
            w199=> c0_n54_w199, 
            w200=> c0_n54_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n54_y
   );           
            
neuron_inst_55: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n55_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n55_w1, 
            w2=> c0_n55_w2, 
            w3=> c0_n55_w3, 
            w4=> c0_n55_w4, 
            w5=> c0_n55_w5, 
            w6=> c0_n55_w6, 
            w7=> c0_n55_w7, 
            w8=> c0_n55_w8, 
            w9=> c0_n55_w9, 
            w10=> c0_n55_w10, 
            w11=> c0_n55_w11, 
            w12=> c0_n55_w12, 
            w13=> c0_n55_w13, 
            w14=> c0_n55_w14, 
            w15=> c0_n55_w15, 
            w16=> c0_n55_w16, 
            w17=> c0_n55_w17, 
            w18=> c0_n55_w18, 
            w19=> c0_n55_w19, 
            w20=> c0_n55_w20, 
            w21=> c0_n55_w21, 
            w22=> c0_n55_w22, 
            w23=> c0_n55_w23, 
            w24=> c0_n55_w24, 
            w25=> c0_n55_w25, 
            w26=> c0_n55_w26, 
            w27=> c0_n55_w27, 
            w28=> c0_n55_w28, 
            w29=> c0_n55_w29, 
            w30=> c0_n55_w30, 
            w31=> c0_n55_w31, 
            w32=> c0_n55_w32, 
            w33=> c0_n55_w33, 
            w34=> c0_n55_w34, 
            w35=> c0_n55_w35, 
            w36=> c0_n55_w36, 
            w37=> c0_n55_w37, 
            w38=> c0_n55_w38, 
            w39=> c0_n55_w39, 
            w40=> c0_n55_w40, 
            w41=> c0_n55_w41, 
            w42=> c0_n55_w42, 
            w43=> c0_n55_w43, 
            w44=> c0_n55_w44, 
            w45=> c0_n55_w45, 
            w46=> c0_n55_w46, 
            w47=> c0_n55_w47, 
            w48=> c0_n55_w48, 
            w49=> c0_n55_w49, 
            w50=> c0_n55_w50, 
            w51=> c0_n55_w51, 
            w52=> c0_n55_w52, 
            w53=> c0_n55_w53, 
            w54=> c0_n55_w54, 
            w55=> c0_n55_w55, 
            w56=> c0_n55_w56, 
            w57=> c0_n55_w57, 
            w58=> c0_n55_w58, 
            w59=> c0_n55_w59, 
            w60=> c0_n55_w60, 
            w61=> c0_n55_w61, 
            w62=> c0_n55_w62, 
            w63=> c0_n55_w63, 
            w64=> c0_n55_w64, 
            w65=> c0_n55_w65, 
            w66=> c0_n55_w66, 
            w67=> c0_n55_w67, 
            w68=> c0_n55_w68, 
            w69=> c0_n55_w69, 
            w70=> c0_n55_w70, 
            w71=> c0_n55_w71, 
            w72=> c0_n55_w72, 
            w73=> c0_n55_w73, 
            w74=> c0_n55_w74, 
            w75=> c0_n55_w75, 
            w76=> c0_n55_w76, 
            w77=> c0_n55_w77, 
            w78=> c0_n55_w78, 
            w79=> c0_n55_w79, 
            w80=> c0_n55_w80, 
            w81=> c0_n55_w81, 
            w82=> c0_n55_w82, 
            w83=> c0_n55_w83, 
            w84=> c0_n55_w84, 
            w85=> c0_n55_w85, 
            w86=> c0_n55_w86, 
            w87=> c0_n55_w87, 
            w88=> c0_n55_w88, 
            w89=> c0_n55_w89, 
            w90=> c0_n55_w90, 
            w91=> c0_n55_w91, 
            w92=> c0_n55_w92, 
            w93=> c0_n55_w93, 
            w94=> c0_n55_w94, 
            w95=> c0_n55_w95, 
            w96=> c0_n55_w96, 
            w97=> c0_n55_w97, 
            w98=> c0_n55_w98, 
            w99=> c0_n55_w99, 
            w100=> c0_n55_w100, 
            w101=> c0_n55_w101, 
            w102=> c0_n55_w102, 
            w103=> c0_n55_w103, 
            w104=> c0_n55_w104, 
            w105=> c0_n55_w105, 
            w106=> c0_n55_w106, 
            w107=> c0_n55_w107, 
            w108=> c0_n55_w108, 
            w109=> c0_n55_w109, 
            w110=> c0_n55_w110, 
            w111=> c0_n55_w111, 
            w112=> c0_n55_w112, 
            w113=> c0_n55_w113, 
            w114=> c0_n55_w114, 
            w115=> c0_n55_w115, 
            w116=> c0_n55_w116, 
            w117=> c0_n55_w117, 
            w118=> c0_n55_w118, 
            w119=> c0_n55_w119, 
            w120=> c0_n55_w120, 
            w121=> c0_n55_w121, 
            w122=> c0_n55_w122, 
            w123=> c0_n55_w123, 
            w124=> c0_n55_w124, 
            w125=> c0_n55_w125, 
            w126=> c0_n55_w126, 
            w127=> c0_n55_w127, 
            w128=> c0_n55_w128, 
            w129=> c0_n55_w129, 
            w130=> c0_n55_w130, 
            w131=> c0_n55_w131, 
            w132=> c0_n55_w132, 
            w133=> c0_n55_w133, 
            w134=> c0_n55_w134, 
            w135=> c0_n55_w135, 
            w136=> c0_n55_w136, 
            w137=> c0_n55_w137, 
            w138=> c0_n55_w138, 
            w139=> c0_n55_w139, 
            w140=> c0_n55_w140, 
            w141=> c0_n55_w141, 
            w142=> c0_n55_w142, 
            w143=> c0_n55_w143, 
            w144=> c0_n55_w144, 
            w145=> c0_n55_w145, 
            w146=> c0_n55_w146, 
            w147=> c0_n55_w147, 
            w148=> c0_n55_w148, 
            w149=> c0_n55_w149, 
            w150=> c0_n55_w150, 
            w151=> c0_n55_w151, 
            w152=> c0_n55_w152, 
            w153=> c0_n55_w153, 
            w154=> c0_n55_w154, 
            w155=> c0_n55_w155, 
            w156=> c0_n55_w156, 
            w157=> c0_n55_w157, 
            w158=> c0_n55_w158, 
            w159=> c0_n55_w159, 
            w160=> c0_n55_w160, 
            w161=> c0_n55_w161, 
            w162=> c0_n55_w162, 
            w163=> c0_n55_w163, 
            w164=> c0_n55_w164, 
            w165=> c0_n55_w165, 
            w166=> c0_n55_w166, 
            w167=> c0_n55_w167, 
            w168=> c0_n55_w168, 
            w169=> c0_n55_w169, 
            w170=> c0_n55_w170, 
            w171=> c0_n55_w171, 
            w172=> c0_n55_w172, 
            w173=> c0_n55_w173, 
            w174=> c0_n55_w174, 
            w175=> c0_n55_w175, 
            w176=> c0_n55_w176, 
            w177=> c0_n55_w177, 
            w178=> c0_n55_w178, 
            w179=> c0_n55_w179, 
            w180=> c0_n55_w180, 
            w181=> c0_n55_w181, 
            w182=> c0_n55_w182, 
            w183=> c0_n55_w183, 
            w184=> c0_n55_w184, 
            w185=> c0_n55_w185, 
            w186=> c0_n55_w186, 
            w187=> c0_n55_w187, 
            w188=> c0_n55_w188, 
            w189=> c0_n55_w189, 
            w190=> c0_n55_w190, 
            w191=> c0_n55_w191, 
            w192=> c0_n55_w192, 
            w193=> c0_n55_w193, 
            w194=> c0_n55_w194, 
            w195=> c0_n55_w195, 
            w196=> c0_n55_w196, 
            w197=> c0_n55_w197, 
            w198=> c0_n55_w198, 
            w199=> c0_n55_w199, 
            w200=> c0_n55_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n55_y
   );           
            
neuron_inst_56: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n56_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n56_w1, 
            w2=> c0_n56_w2, 
            w3=> c0_n56_w3, 
            w4=> c0_n56_w4, 
            w5=> c0_n56_w5, 
            w6=> c0_n56_w6, 
            w7=> c0_n56_w7, 
            w8=> c0_n56_w8, 
            w9=> c0_n56_w9, 
            w10=> c0_n56_w10, 
            w11=> c0_n56_w11, 
            w12=> c0_n56_w12, 
            w13=> c0_n56_w13, 
            w14=> c0_n56_w14, 
            w15=> c0_n56_w15, 
            w16=> c0_n56_w16, 
            w17=> c0_n56_w17, 
            w18=> c0_n56_w18, 
            w19=> c0_n56_w19, 
            w20=> c0_n56_w20, 
            w21=> c0_n56_w21, 
            w22=> c0_n56_w22, 
            w23=> c0_n56_w23, 
            w24=> c0_n56_w24, 
            w25=> c0_n56_w25, 
            w26=> c0_n56_w26, 
            w27=> c0_n56_w27, 
            w28=> c0_n56_w28, 
            w29=> c0_n56_w29, 
            w30=> c0_n56_w30, 
            w31=> c0_n56_w31, 
            w32=> c0_n56_w32, 
            w33=> c0_n56_w33, 
            w34=> c0_n56_w34, 
            w35=> c0_n56_w35, 
            w36=> c0_n56_w36, 
            w37=> c0_n56_w37, 
            w38=> c0_n56_w38, 
            w39=> c0_n56_w39, 
            w40=> c0_n56_w40, 
            w41=> c0_n56_w41, 
            w42=> c0_n56_w42, 
            w43=> c0_n56_w43, 
            w44=> c0_n56_w44, 
            w45=> c0_n56_w45, 
            w46=> c0_n56_w46, 
            w47=> c0_n56_w47, 
            w48=> c0_n56_w48, 
            w49=> c0_n56_w49, 
            w50=> c0_n56_w50, 
            w51=> c0_n56_w51, 
            w52=> c0_n56_w52, 
            w53=> c0_n56_w53, 
            w54=> c0_n56_w54, 
            w55=> c0_n56_w55, 
            w56=> c0_n56_w56, 
            w57=> c0_n56_w57, 
            w58=> c0_n56_w58, 
            w59=> c0_n56_w59, 
            w60=> c0_n56_w60, 
            w61=> c0_n56_w61, 
            w62=> c0_n56_w62, 
            w63=> c0_n56_w63, 
            w64=> c0_n56_w64, 
            w65=> c0_n56_w65, 
            w66=> c0_n56_w66, 
            w67=> c0_n56_w67, 
            w68=> c0_n56_w68, 
            w69=> c0_n56_w69, 
            w70=> c0_n56_w70, 
            w71=> c0_n56_w71, 
            w72=> c0_n56_w72, 
            w73=> c0_n56_w73, 
            w74=> c0_n56_w74, 
            w75=> c0_n56_w75, 
            w76=> c0_n56_w76, 
            w77=> c0_n56_w77, 
            w78=> c0_n56_w78, 
            w79=> c0_n56_w79, 
            w80=> c0_n56_w80, 
            w81=> c0_n56_w81, 
            w82=> c0_n56_w82, 
            w83=> c0_n56_w83, 
            w84=> c0_n56_w84, 
            w85=> c0_n56_w85, 
            w86=> c0_n56_w86, 
            w87=> c0_n56_w87, 
            w88=> c0_n56_w88, 
            w89=> c0_n56_w89, 
            w90=> c0_n56_w90, 
            w91=> c0_n56_w91, 
            w92=> c0_n56_w92, 
            w93=> c0_n56_w93, 
            w94=> c0_n56_w94, 
            w95=> c0_n56_w95, 
            w96=> c0_n56_w96, 
            w97=> c0_n56_w97, 
            w98=> c0_n56_w98, 
            w99=> c0_n56_w99, 
            w100=> c0_n56_w100, 
            w101=> c0_n56_w101, 
            w102=> c0_n56_w102, 
            w103=> c0_n56_w103, 
            w104=> c0_n56_w104, 
            w105=> c0_n56_w105, 
            w106=> c0_n56_w106, 
            w107=> c0_n56_w107, 
            w108=> c0_n56_w108, 
            w109=> c0_n56_w109, 
            w110=> c0_n56_w110, 
            w111=> c0_n56_w111, 
            w112=> c0_n56_w112, 
            w113=> c0_n56_w113, 
            w114=> c0_n56_w114, 
            w115=> c0_n56_w115, 
            w116=> c0_n56_w116, 
            w117=> c0_n56_w117, 
            w118=> c0_n56_w118, 
            w119=> c0_n56_w119, 
            w120=> c0_n56_w120, 
            w121=> c0_n56_w121, 
            w122=> c0_n56_w122, 
            w123=> c0_n56_w123, 
            w124=> c0_n56_w124, 
            w125=> c0_n56_w125, 
            w126=> c0_n56_w126, 
            w127=> c0_n56_w127, 
            w128=> c0_n56_w128, 
            w129=> c0_n56_w129, 
            w130=> c0_n56_w130, 
            w131=> c0_n56_w131, 
            w132=> c0_n56_w132, 
            w133=> c0_n56_w133, 
            w134=> c0_n56_w134, 
            w135=> c0_n56_w135, 
            w136=> c0_n56_w136, 
            w137=> c0_n56_w137, 
            w138=> c0_n56_w138, 
            w139=> c0_n56_w139, 
            w140=> c0_n56_w140, 
            w141=> c0_n56_w141, 
            w142=> c0_n56_w142, 
            w143=> c0_n56_w143, 
            w144=> c0_n56_w144, 
            w145=> c0_n56_w145, 
            w146=> c0_n56_w146, 
            w147=> c0_n56_w147, 
            w148=> c0_n56_w148, 
            w149=> c0_n56_w149, 
            w150=> c0_n56_w150, 
            w151=> c0_n56_w151, 
            w152=> c0_n56_w152, 
            w153=> c0_n56_w153, 
            w154=> c0_n56_w154, 
            w155=> c0_n56_w155, 
            w156=> c0_n56_w156, 
            w157=> c0_n56_w157, 
            w158=> c0_n56_w158, 
            w159=> c0_n56_w159, 
            w160=> c0_n56_w160, 
            w161=> c0_n56_w161, 
            w162=> c0_n56_w162, 
            w163=> c0_n56_w163, 
            w164=> c0_n56_w164, 
            w165=> c0_n56_w165, 
            w166=> c0_n56_w166, 
            w167=> c0_n56_w167, 
            w168=> c0_n56_w168, 
            w169=> c0_n56_w169, 
            w170=> c0_n56_w170, 
            w171=> c0_n56_w171, 
            w172=> c0_n56_w172, 
            w173=> c0_n56_w173, 
            w174=> c0_n56_w174, 
            w175=> c0_n56_w175, 
            w176=> c0_n56_w176, 
            w177=> c0_n56_w177, 
            w178=> c0_n56_w178, 
            w179=> c0_n56_w179, 
            w180=> c0_n56_w180, 
            w181=> c0_n56_w181, 
            w182=> c0_n56_w182, 
            w183=> c0_n56_w183, 
            w184=> c0_n56_w184, 
            w185=> c0_n56_w185, 
            w186=> c0_n56_w186, 
            w187=> c0_n56_w187, 
            w188=> c0_n56_w188, 
            w189=> c0_n56_w189, 
            w190=> c0_n56_w190, 
            w191=> c0_n56_w191, 
            w192=> c0_n56_w192, 
            w193=> c0_n56_w193, 
            w194=> c0_n56_w194, 
            w195=> c0_n56_w195, 
            w196=> c0_n56_w196, 
            w197=> c0_n56_w197, 
            w198=> c0_n56_w198, 
            w199=> c0_n56_w199, 
            w200=> c0_n56_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n56_y
   );           
            
neuron_inst_57: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n57_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n57_w1, 
            w2=> c0_n57_w2, 
            w3=> c0_n57_w3, 
            w4=> c0_n57_w4, 
            w5=> c0_n57_w5, 
            w6=> c0_n57_w6, 
            w7=> c0_n57_w7, 
            w8=> c0_n57_w8, 
            w9=> c0_n57_w9, 
            w10=> c0_n57_w10, 
            w11=> c0_n57_w11, 
            w12=> c0_n57_w12, 
            w13=> c0_n57_w13, 
            w14=> c0_n57_w14, 
            w15=> c0_n57_w15, 
            w16=> c0_n57_w16, 
            w17=> c0_n57_w17, 
            w18=> c0_n57_w18, 
            w19=> c0_n57_w19, 
            w20=> c0_n57_w20, 
            w21=> c0_n57_w21, 
            w22=> c0_n57_w22, 
            w23=> c0_n57_w23, 
            w24=> c0_n57_w24, 
            w25=> c0_n57_w25, 
            w26=> c0_n57_w26, 
            w27=> c0_n57_w27, 
            w28=> c0_n57_w28, 
            w29=> c0_n57_w29, 
            w30=> c0_n57_w30, 
            w31=> c0_n57_w31, 
            w32=> c0_n57_w32, 
            w33=> c0_n57_w33, 
            w34=> c0_n57_w34, 
            w35=> c0_n57_w35, 
            w36=> c0_n57_w36, 
            w37=> c0_n57_w37, 
            w38=> c0_n57_w38, 
            w39=> c0_n57_w39, 
            w40=> c0_n57_w40, 
            w41=> c0_n57_w41, 
            w42=> c0_n57_w42, 
            w43=> c0_n57_w43, 
            w44=> c0_n57_w44, 
            w45=> c0_n57_w45, 
            w46=> c0_n57_w46, 
            w47=> c0_n57_w47, 
            w48=> c0_n57_w48, 
            w49=> c0_n57_w49, 
            w50=> c0_n57_w50, 
            w51=> c0_n57_w51, 
            w52=> c0_n57_w52, 
            w53=> c0_n57_w53, 
            w54=> c0_n57_w54, 
            w55=> c0_n57_w55, 
            w56=> c0_n57_w56, 
            w57=> c0_n57_w57, 
            w58=> c0_n57_w58, 
            w59=> c0_n57_w59, 
            w60=> c0_n57_w60, 
            w61=> c0_n57_w61, 
            w62=> c0_n57_w62, 
            w63=> c0_n57_w63, 
            w64=> c0_n57_w64, 
            w65=> c0_n57_w65, 
            w66=> c0_n57_w66, 
            w67=> c0_n57_w67, 
            w68=> c0_n57_w68, 
            w69=> c0_n57_w69, 
            w70=> c0_n57_w70, 
            w71=> c0_n57_w71, 
            w72=> c0_n57_w72, 
            w73=> c0_n57_w73, 
            w74=> c0_n57_w74, 
            w75=> c0_n57_w75, 
            w76=> c0_n57_w76, 
            w77=> c0_n57_w77, 
            w78=> c0_n57_w78, 
            w79=> c0_n57_w79, 
            w80=> c0_n57_w80, 
            w81=> c0_n57_w81, 
            w82=> c0_n57_w82, 
            w83=> c0_n57_w83, 
            w84=> c0_n57_w84, 
            w85=> c0_n57_w85, 
            w86=> c0_n57_w86, 
            w87=> c0_n57_w87, 
            w88=> c0_n57_w88, 
            w89=> c0_n57_w89, 
            w90=> c0_n57_w90, 
            w91=> c0_n57_w91, 
            w92=> c0_n57_w92, 
            w93=> c0_n57_w93, 
            w94=> c0_n57_w94, 
            w95=> c0_n57_w95, 
            w96=> c0_n57_w96, 
            w97=> c0_n57_w97, 
            w98=> c0_n57_w98, 
            w99=> c0_n57_w99, 
            w100=> c0_n57_w100, 
            w101=> c0_n57_w101, 
            w102=> c0_n57_w102, 
            w103=> c0_n57_w103, 
            w104=> c0_n57_w104, 
            w105=> c0_n57_w105, 
            w106=> c0_n57_w106, 
            w107=> c0_n57_w107, 
            w108=> c0_n57_w108, 
            w109=> c0_n57_w109, 
            w110=> c0_n57_w110, 
            w111=> c0_n57_w111, 
            w112=> c0_n57_w112, 
            w113=> c0_n57_w113, 
            w114=> c0_n57_w114, 
            w115=> c0_n57_w115, 
            w116=> c0_n57_w116, 
            w117=> c0_n57_w117, 
            w118=> c0_n57_w118, 
            w119=> c0_n57_w119, 
            w120=> c0_n57_w120, 
            w121=> c0_n57_w121, 
            w122=> c0_n57_w122, 
            w123=> c0_n57_w123, 
            w124=> c0_n57_w124, 
            w125=> c0_n57_w125, 
            w126=> c0_n57_w126, 
            w127=> c0_n57_w127, 
            w128=> c0_n57_w128, 
            w129=> c0_n57_w129, 
            w130=> c0_n57_w130, 
            w131=> c0_n57_w131, 
            w132=> c0_n57_w132, 
            w133=> c0_n57_w133, 
            w134=> c0_n57_w134, 
            w135=> c0_n57_w135, 
            w136=> c0_n57_w136, 
            w137=> c0_n57_w137, 
            w138=> c0_n57_w138, 
            w139=> c0_n57_w139, 
            w140=> c0_n57_w140, 
            w141=> c0_n57_w141, 
            w142=> c0_n57_w142, 
            w143=> c0_n57_w143, 
            w144=> c0_n57_w144, 
            w145=> c0_n57_w145, 
            w146=> c0_n57_w146, 
            w147=> c0_n57_w147, 
            w148=> c0_n57_w148, 
            w149=> c0_n57_w149, 
            w150=> c0_n57_w150, 
            w151=> c0_n57_w151, 
            w152=> c0_n57_w152, 
            w153=> c0_n57_w153, 
            w154=> c0_n57_w154, 
            w155=> c0_n57_w155, 
            w156=> c0_n57_w156, 
            w157=> c0_n57_w157, 
            w158=> c0_n57_w158, 
            w159=> c0_n57_w159, 
            w160=> c0_n57_w160, 
            w161=> c0_n57_w161, 
            w162=> c0_n57_w162, 
            w163=> c0_n57_w163, 
            w164=> c0_n57_w164, 
            w165=> c0_n57_w165, 
            w166=> c0_n57_w166, 
            w167=> c0_n57_w167, 
            w168=> c0_n57_w168, 
            w169=> c0_n57_w169, 
            w170=> c0_n57_w170, 
            w171=> c0_n57_w171, 
            w172=> c0_n57_w172, 
            w173=> c0_n57_w173, 
            w174=> c0_n57_w174, 
            w175=> c0_n57_w175, 
            w176=> c0_n57_w176, 
            w177=> c0_n57_w177, 
            w178=> c0_n57_w178, 
            w179=> c0_n57_w179, 
            w180=> c0_n57_w180, 
            w181=> c0_n57_w181, 
            w182=> c0_n57_w182, 
            w183=> c0_n57_w183, 
            w184=> c0_n57_w184, 
            w185=> c0_n57_w185, 
            w186=> c0_n57_w186, 
            w187=> c0_n57_w187, 
            w188=> c0_n57_w188, 
            w189=> c0_n57_w189, 
            w190=> c0_n57_w190, 
            w191=> c0_n57_w191, 
            w192=> c0_n57_w192, 
            w193=> c0_n57_w193, 
            w194=> c0_n57_w194, 
            w195=> c0_n57_w195, 
            w196=> c0_n57_w196, 
            w197=> c0_n57_w197, 
            w198=> c0_n57_w198, 
            w199=> c0_n57_w199, 
            w200=> c0_n57_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n57_y
   );           
            
neuron_inst_58: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n58_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n58_w1, 
            w2=> c0_n58_w2, 
            w3=> c0_n58_w3, 
            w4=> c0_n58_w4, 
            w5=> c0_n58_w5, 
            w6=> c0_n58_w6, 
            w7=> c0_n58_w7, 
            w8=> c0_n58_w8, 
            w9=> c0_n58_w9, 
            w10=> c0_n58_w10, 
            w11=> c0_n58_w11, 
            w12=> c0_n58_w12, 
            w13=> c0_n58_w13, 
            w14=> c0_n58_w14, 
            w15=> c0_n58_w15, 
            w16=> c0_n58_w16, 
            w17=> c0_n58_w17, 
            w18=> c0_n58_w18, 
            w19=> c0_n58_w19, 
            w20=> c0_n58_w20, 
            w21=> c0_n58_w21, 
            w22=> c0_n58_w22, 
            w23=> c0_n58_w23, 
            w24=> c0_n58_w24, 
            w25=> c0_n58_w25, 
            w26=> c0_n58_w26, 
            w27=> c0_n58_w27, 
            w28=> c0_n58_w28, 
            w29=> c0_n58_w29, 
            w30=> c0_n58_w30, 
            w31=> c0_n58_w31, 
            w32=> c0_n58_w32, 
            w33=> c0_n58_w33, 
            w34=> c0_n58_w34, 
            w35=> c0_n58_w35, 
            w36=> c0_n58_w36, 
            w37=> c0_n58_w37, 
            w38=> c0_n58_w38, 
            w39=> c0_n58_w39, 
            w40=> c0_n58_w40, 
            w41=> c0_n58_w41, 
            w42=> c0_n58_w42, 
            w43=> c0_n58_w43, 
            w44=> c0_n58_w44, 
            w45=> c0_n58_w45, 
            w46=> c0_n58_w46, 
            w47=> c0_n58_w47, 
            w48=> c0_n58_w48, 
            w49=> c0_n58_w49, 
            w50=> c0_n58_w50, 
            w51=> c0_n58_w51, 
            w52=> c0_n58_w52, 
            w53=> c0_n58_w53, 
            w54=> c0_n58_w54, 
            w55=> c0_n58_w55, 
            w56=> c0_n58_w56, 
            w57=> c0_n58_w57, 
            w58=> c0_n58_w58, 
            w59=> c0_n58_w59, 
            w60=> c0_n58_w60, 
            w61=> c0_n58_w61, 
            w62=> c0_n58_w62, 
            w63=> c0_n58_w63, 
            w64=> c0_n58_w64, 
            w65=> c0_n58_w65, 
            w66=> c0_n58_w66, 
            w67=> c0_n58_w67, 
            w68=> c0_n58_w68, 
            w69=> c0_n58_w69, 
            w70=> c0_n58_w70, 
            w71=> c0_n58_w71, 
            w72=> c0_n58_w72, 
            w73=> c0_n58_w73, 
            w74=> c0_n58_w74, 
            w75=> c0_n58_w75, 
            w76=> c0_n58_w76, 
            w77=> c0_n58_w77, 
            w78=> c0_n58_w78, 
            w79=> c0_n58_w79, 
            w80=> c0_n58_w80, 
            w81=> c0_n58_w81, 
            w82=> c0_n58_w82, 
            w83=> c0_n58_w83, 
            w84=> c0_n58_w84, 
            w85=> c0_n58_w85, 
            w86=> c0_n58_w86, 
            w87=> c0_n58_w87, 
            w88=> c0_n58_w88, 
            w89=> c0_n58_w89, 
            w90=> c0_n58_w90, 
            w91=> c0_n58_w91, 
            w92=> c0_n58_w92, 
            w93=> c0_n58_w93, 
            w94=> c0_n58_w94, 
            w95=> c0_n58_w95, 
            w96=> c0_n58_w96, 
            w97=> c0_n58_w97, 
            w98=> c0_n58_w98, 
            w99=> c0_n58_w99, 
            w100=> c0_n58_w100, 
            w101=> c0_n58_w101, 
            w102=> c0_n58_w102, 
            w103=> c0_n58_w103, 
            w104=> c0_n58_w104, 
            w105=> c0_n58_w105, 
            w106=> c0_n58_w106, 
            w107=> c0_n58_w107, 
            w108=> c0_n58_w108, 
            w109=> c0_n58_w109, 
            w110=> c0_n58_w110, 
            w111=> c0_n58_w111, 
            w112=> c0_n58_w112, 
            w113=> c0_n58_w113, 
            w114=> c0_n58_w114, 
            w115=> c0_n58_w115, 
            w116=> c0_n58_w116, 
            w117=> c0_n58_w117, 
            w118=> c0_n58_w118, 
            w119=> c0_n58_w119, 
            w120=> c0_n58_w120, 
            w121=> c0_n58_w121, 
            w122=> c0_n58_w122, 
            w123=> c0_n58_w123, 
            w124=> c0_n58_w124, 
            w125=> c0_n58_w125, 
            w126=> c0_n58_w126, 
            w127=> c0_n58_w127, 
            w128=> c0_n58_w128, 
            w129=> c0_n58_w129, 
            w130=> c0_n58_w130, 
            w131=> c0_n58_w131, 
            w132=> c0_n58_w132, 
            w133=> c0_n58_w133, 
            w134=> c0_n58_w134, 
            w135=> c0_n58_w135, 
            w136=> c0_n58_w136, 
            w137=> c0_n58_w137, 
            w138=> c0_n58_w138, 
            w139=> c0_n58_w139, 
            w140=> c0_n58_w140, 
            w141=> c0_n58_w141, 
            w142=> c0_n58_w142, 
            w143=> c0_n58_w143, 
            w144=> c0_n58_w144, 
            w145=> c0_n58_w145, 
            w146=> c0_n58_w146, 
            w147=> c0_n58_w147, 
            w148=> c0_n58_w148, 
            w149=> c0_n58_w149, 
            w150=> c0_n58_w150, 
            w151=> c0_n58_w151, 
            w152=> c0_n58_w152, 
            w153=> c0_n58_w153, 
            w154=> c0_n58_w154, 
            w155=> c0_n58_w155, 
            w156=> c0_n58_w156, 
            w157=> c0_n58_w157, 
            w158=> c0_n58_w158, 
            w159=> c0_n58_w159, 
            w160=> c0_n58_w160, 
            w161=> c0_n58_w161, 
            w162=> c0_n58_w162, 
            w163=> c0_n58_w163, 
            w164=> c0_n58_w164, 
            w165=> c0_n58_w165, 
            w166=> c0_n58_w166, 
            w167=> c0_n58_w167, 
            w168=> c0_n58_w168, 
            w169=> c0_n58_w169, 
            w170=> c0_n58_w170, 
            w171=> c0_n58_w171, 
            w172=> c0_n58_w172, 
            w173=> c0_n58_w173, 
            w174=> c0_n58_w174, 
            w175=> c0_n58_w175, 
            w176=> c0_n58_w176, 
            w177=> c0_n58_w177, 
            w178=> c0_n58_w178, 
            w179=> c0_n58_w179, 
            w180=> c0_n58_w180, 
            w181=> c0_n58_w181, 
            w182=> c0_n58_w182, 
            w183=> c0_n58_w183, 
            w184=> c0_n58_w184, 
            w185=> c0_n58_w185, 
            w186=> c0_n58_w186, 
            w187=> c0_n58_w187, 
            w188=> c0_n58_w188, 
            w189=> c0_n58_w189, 
            w190=> c0_n58_w190, 
            w191=> c0_n58_w191, 
            w192=> c0_n58_w192, 
            w193=> c0_n58_w193, 
            w194=> c0_n58_w194, 
            w195=> c0_n58_w195, 
            w196=> c0_n58_w196, 
            w197=> c0_n58_w197, 
            w198=> c0_n58_w198, 
            w199=> c0_n58_w199, 
            w200=> c0_n58_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n58_y
   );           
            
neuron_inst_59: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n59_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n59_w1, 
            w2=> c0_n59_w2, 
            w3=> c0_n59_w3, 
            w4=> c0_n59_w4, 
            w5=> c0_n59_w5, 
            w6=> c0_n59_w6, 
            w7=> c0_n59_w7, 
            w8=> c0_n59_w8, 
            w9=> c0_n59_w9, 
            w10=> c0_n59_w10, 
            w11=> c0_n59_w11, 
            w12=> c0_n59_w12, 
            w13=> c0_n59_w13, 
            w14=> c0_n59_w14, 
            w15=> c0_n59_w15, 
            w16=> c0_n59_w16, 
            w17=> c0_n59_w17, 
            w18=> c0_n59_w18, 
            w19=> c0_n59_w19, 
            w20=> c0_n59_w20, 
            w21=> c0_n59_w21, 
            w22=> c0_n59_w22, 
            w23=> c0_n59_w23, 
            w24=> c0_n59_w24, 
            w25=> c0_n59_w25, 
            w26=> c0_n59_w26, 
            w27=> c0_n59_w27, 
            w28=> c0_n59_w28, 
            w29=> c0_n59_w29, 
            w30=> c0_n59_w30, 
            w31=> c0_n59_w31, 
            w32=> c0_n59_w32, 
            w33=> c0_n59_w33, 
            w34=> c0_n59_w34, 
            w35=> c0_n59_w35, 
            w36=> c0_n59_w36, 
            w37=> c0_n59_w37, 
            w38=> c0_n59_w38, 
            w39=> c0_n59_w39, 
            w40=> c0_n59_w40, 
            w41=> c0_n59_w41, 
            w42=> c0_n59_w42, 
            w43=> c0_n59_w43, 
            w44=> c0_n59_w44, 
            w45=> c0_n59_w45, 
            w46=> c0_n59_w46, 
            w47=> c0_n59_w47, 
            w48=> c0_n59_w48, 
            w49=> c0_n59_w49, 
            w50=> c0_n59_w50, 
            w51=> c0_n59_w51, 
            w52=> c0_n59_w52, 
            w53=> c0_n59_w53, 
            w54=> c0_n59_w54, 
            w55=> c0_n59_w55, 
            w56=> c0_n59_w56, 
            w57=> c0_n59_w57, 
            w58=> c0_n59_w58, 
            w59=> c0_n59_w59, 
            w60=> c0_n59_w60, 
            w61=> c0_n59_w61, 
            w62=> c0_n59_w62, 
            w63=> c0_n59_w63, 
            w64=> c0_n59_w64, 
            w65=> c0_n59_w65, 
            w66=> c0_n59_w66, 
            w67=> c0_n59_w67, 
            w68=> c0_n59_w68, 
            w69=> c0_n59_w69, 
            w70=> c0_n59_w70, 
            w71=> c0_n59_w71, 
            w72=> c0_n59_w72, 
            w73=> c0_n59_w73, 
            w74=> c0_n59_w74, 
            w75=> c0_n59_w75, 
            w76=> c0_n59_w76, 
            w77=> c0_n59_w77, 
            w78=> c0_n59_w78, 
            w79=> c0_n59_w79, 
            w80=> c0_n59_w80, 
            w81=> c0_n59_w81, 
            w82=> c0_n59_w82, 
            w83=> c0_n59_w83, 
            w84=> c0_n59_w84, 
            w85=> c0_n59_w85, 
            w86=> c0_n59_w86, 
            w87=> c0_n59_w87, 
            w88=> c0_n59_w88, 
            w89=> c0_n59_w89, 
            w90=> c0_n59_w90, 
            w91=> c0_n59_w91, 
            w92=> c0_n59_w92, 
            w93=> c0_n59_w93, 
            w94=> c0_n59_w94, 
            w95=> c0_n59_w95, 
            w96=> c0_n59_w96, 
            w97=> c0_n59_w97, 
            w98=> c0_n59_w98, 
            w99=> c0_n59_w99, 
            w100=> c0_n59_w100, 
            w101=> c0_n59_w101, 
            w102=> c0_n59_w102, 
            w103=> c0_n59_w103, 
            w104=> c0_n59_w104, 
            w105=> c0_n59_w105, 
            w106=> c0_n59_w106, 
            w107=> c0_n59_w107, 
            w108=> c0_n59_w108, 
            w109=> c0_n59_w109, 
            w110=> c0_n59_w110, 
            w111=> c0_n59_w111, 
            w112=> c0_n59_w112, 
            w113=> c0_n59_w113, 
            w114=> c0_n59_w114, 
            w115=> c0_n59_w115, 
            w116=> c0_n59_w116, 
            w117=> c0_n59_w117, 
            w118=> c0_n59_w118, 
            w119=> c0_n59_w119, 
            w120=> c0_n59_w120, 
            w121=> c0_n59_w121, 
            w122=> c0_n59_w122, 
            w123=> c0_n59_w123, 
            w124=> c0_n59_w124, 
            w125=> c0_n59_w125, 
            w126=> c0_n59_w126, 
            w127=> c0_n59_w127, 
            w128=> c0_n59_w128, 
            w129=> c0_n59_w129, 
            w130=> c0_n59_w130, 
            w131=> c0_n59_w131, 
            w132=> c0_n59_w132, 
            w133=> c0_n59_w133, 
            w134=> c0_n59_w134, 
            w135=> c0_n59_w135, 
            w136=> c0_n59_w136, 
            w137=> c0_n59_w137, 
            w138=> c0_n59_w138, 
            w139=> c0_n59_w139, 
            w140=> c0_n59_w140, 
            w141=> c0_n59_w141, 
            w142=> c0_n59_w142, 
            w143=> c0_n59_w143, 
            w144=> c0_n59_w144, 
            w145=> c0_n59_w145, 
            w146=> c0_n59_w146, 
            w147=> c0_n59_w147, 
            w148=> c0_n59_w148, 
            w149=> c0_n59_w149, 
            w150=> c0_n59_w150, 
            w151=> c0_n59_w151, 
            w152=> c0_n59_w152, 
            w153=> c0_n59_w153, 
            w154=> c0_n59_w154, 
            w155=> c0_n59_w155, 
            w156=> c0_n59_w156, 
            w157=> c0_n59_w157, 
            w158=> c0_n59_w158, 
            w159=> c0_n59_w159, 
            w160=> c0_n59_w160, 
            w161=> c0_n59_w161, 
            w162=> c0_n59_w162, 
            w163=> c0_n59_w163, 
            w164=> c0_n59_w164, 
            w165=> c0_n59_w165, 
            w166=> c0_n59_w166, 
            w167=> c0_n59_w167, 
            w168=> c0_n59_w168, 
            w169=> c0_n59_w169, 
            w170=> c0_n59_w170, 
            w171=> c0_n59_w171, 
            w172=> c0_n59_w172, 
            w173=> c0_n59_w173, 
            w174=> c0_n59_w174, 
            w175=> c0_n59_w175, 
            w176=> c0_n59_w176, 
            w177=> c0_n59_w177, 
            w178=> c0_n59_w178, 
            w179=> c0_n59_w179, 
            w180=> c0_n59_w180, 
            w181=> c0_n59_w181, 
            w182=> c0_n59_w182, 
            w183=> c0_n59_w183, 
            w184=> c0_n59_w184, 
            w185=> c0_n59_w185, 
            w186=> c0_n59_w186, 
            w187=> c0_n59_w187, 
            w188=> c0_n59_w188, 
            w189=> c0_n59_w189, 
            w190=> c0_n59_w190, 
            w191=> c0_n59_w191, 
            w192=> c0_n59_w192, 
            w193=> c0_n59_w193, 
            w194=> c0_n59_w194, 
            w195=> c0_n59_w195, 
            w196=> c0_n59_w196, 
            w197=> c0_n59_w197, 
            w198=> c0_n59_w198, 
            w199=> c0_n59_w199, 
            w200=> c0_n59_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n59_y
   );           
            
neuron_inst_60: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n60_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n60_w1, 
            w2=> c0_n60_w2, 
            w3=> c0_n60_w3, 
            w4=> c0_n60_w4, 
            w5=> c0_n60_w5, 
            w6=> c0_n60_w6, 
            w7=> c0_n60_w7, 
            w8=> c0_n60_w8, 
            w9=> c0_n60_w9, 
            w10=> c0_n60_w10, 
            w11=> c0_n60_w11, 
            w12=> c0_n60_w12, 
            w13=> c0_n60_w13, 
            w14=> c0_n60_w14, 
            w15=> c0_n60_w15, 
            w16=> c0_n60_w16, 
            w17=> c0_n60_w17, 
            w18=> c0_n60_w18, 
            w19=> c0_n60_w19, 
            w20=> c0_n60_w20, 
            w21=> c0_n60_w21, 
            w22=> c0_n60_w22, 
            w23=> c0_n60_w23, 
            w24=> c0_n60_w24, 
            w25=> c0_n60_w25, 
            w26=> c0_n60_w26, 
            w27=> c0_n60_w27, 
            w28=> c0_n60_w28, 
            w29=> c0_n60_w29, 
            w30=> c0_n60_w30, 
            w31=> c0_n60_w31, 
            w32=> c0_n60_w32, 
            w33=> c0_n60_w33, 
            w34=> c0_n60_w34, 
            w35=> c0_n60_w35, 
            w36=> c0_n60_w36, 
            w37=> c0_n60_w37, 
            w38=> c0_n60_w38, 
            w39=> c0_n60_w39, 
            w40=> c0_n60_w40, 
            w41=> c0_n60_w41, 
            w42=> c0_n60_w42, 
            w43=> c0_n60_w43, 
            w44=> c0_n60_w44, 
            w45=> c0_n60_w45, 
            w46=> c0_n60_w46, 
            w47=> c0_n60_w47, 
            w48=> c0_n60_w48, 
            w49=> c0_n60_w49, 
            w50=> c0_n60_w50, 
            w51=> c0_n60_w51, 
            w52=> c0_n60_w52, 
            w53=> c0_n60_w53, 
            w54=> c0_n60_w54, 
            w55=> c0_n60_w55, 
            w56=> c0_n60_w56, 
            w57=> c0_n60_w57, 
            w58=> c0_n60_w58, 
            w59=> c0_n60_w59, 
            w60=> c0_n60_w60, 
            w61=> c0_n60_w61, 
            w62=> c0_n60_w62, 
            w63=> c0_n60_w63, 
            w64=> c0_n60_w64, 
            w65=> c0_n60_w65, 
            w66=> c0_n60_w66, 
            w67=> c0_n60_w67, 
            w68=> c0_n60_w68, 
            w69=> c0_n60_w69, 
            w70=> c0_n60_w70, 
            w71=> c0_n60_w71, 
            w72=> c0_n60_w72, 
            w73=> c0_n60_w73, 
            w74=> c0_n60_w74, 
            w75=> c0_n60_w75, 
            w76=> c0_n60_w76, 
            w77=> c0_n60_w77, 
            w78=> c0_n60_w78, 
            w79=> c0_n60_w79, 
            w80=> c0_n60_w80, 
            w81=> c0_n60_w81, 
            w82=> c0_n60_w82, 
            w83=> c0_n60_w83, 
            w84=> c0_n60_w84, 
            w85=> c0_n60_w85, 
            w86=> c0_n60_w86, 
            w87=> c0_n60_w87, 
            w88=> c0_n60_w88, 
            w89=> c0_n60_w89, 
            w90=> c0_n60_w90, 
            w91=> c0_n60_w91, 
            w92=> c0_n60_w92, 
            w93=> c0_n60_w93, 
            w94=> c0_n60_w94, 
            w95=> c0_n60_w95, 
            w96=> c0_n60_w96, 
            w97=> c0_n60_w97, 
            w98=> c0_n60_w98, 
            w99=> c0_n60_w99, 
            w100=> c0_n60_w100, 
            w101=> c0_n60_w101, 
            w102=> c0_n60_w102, 
            w103=> c0_n60_w103, 
            w104=> c0_n60_w104, 
            w105=> c0_n60_w105, 
            w106=> c0_n60_w106, 
            w107=> c0_n60_w107, 
            w108=> c0_n60_w108, 
            w109=> c0_n60_w109, 
            w110=> c0_n60_w110, 
            w111=> c0_n60_w111, 
            w112=> c0_n60_w112, 
            w113=> c0_n60_w113, 
            w114=> c0_n60_w114, 
            w115=> c0_n60_w115, 
            w116=> c0_n60_w116, 
            w117=> c0_n60_w117, 
            w118=> c0_n60_w118, 
            w119=> c0_n60_w119, 
            w120=> c0_n60_w120, 
            w121=> c0_n60_w121, 
            w122=> c0_n60_w122, 
            w123=> c0_n60_w123, 
            w124=> c0_n60_w124, 
            w125=> c0_n60_w125, 
            w126=> c0_n60_w126, 
            w127=> c0_n60_w127, 
            w128=> c0_n60_w128, 
            w129=> c0_n60_w129, 
            w130=> c0_n60_w130, 
            w131=> c0_n60_w131, 
            w132=> c0_n60_w132, 
            w133=> c0_n60_w133, 
            w134=> c0_n60_w134, 
            w135=> c0_n60_w135, 
            w136=> c0_n60_w136, 
            w137=> c0_n60_w137, 
            w138=> c0_n60_w138, 
            w139=> c0_n60_w139, 
            w140=> c0_n60_w140, 
            w141=> c0_n60_w141, 
            w142=> c0_n60_w142, 
            w143=> c0_n60_w143, 
            w144=> c0_n60_w144, 
            w145=> c0_n60_w145, 
            w146=> c0_n60_w146, 
            w147=> c0_n60_w147, 
            w148=> c0_n60_w148, 
            w149=> c0_n60_w149, 
            w150=> c0_n60_w150, 
            w151=> c0_n60_w151, 
            w152=> c0_n60_w152, 
            w153=> c0_n60_w153, 
            w154=> c0_n60_w154, 
            w155=> c0_n60_w155, 
            w156=> c0_n60_w156, 
            w157=> c0_n60_w157, 
            w158=> c0_n60_w158, 
            w159=> c0_n60_w159, 
            w160=> c0_n60_w160, 
            w161=> c0_n60_w161, 
            w162=> c0_n60_w162, 
            w163=> c0_n60_w163, 
            w164=> c0_n60_w164, 
            w165=> c0_n60_w165, 
            w166=> c0_n60_w166, 
            w167=> c0_n60_w167, 
            w168=> c0_n60_w168, 
            w169=> c0_n60_w169, 
            w170=> c0_n60_w170, 
            w171=> c0_n60_w171, 
            w172=> c0_n60_w172, 
            w173=> c0_n60_w173, 
            w174=> c0_n60_w174, 
            w175=> c0_n60_w175, 
            w176=> c0_n60_w176, 
            w177=> c0_n60_w177, 
            w178=> c0_n60_w178, 
            w179=> c0_n60_w179, 
            w180=> c0_n60_w180, 
            w181=> c0_n60_w181, 
            w182=> c0_n60_w182, 
            w183=> c0_n60_w183, 
            w184=> c0_n60_w184, 
            w185=> c0_n60_w185, 
            w186=> c0_n60_w186, 
            w187=> c0_n60_w187, 
            w188=> c0_n60_w188, 
            w189=> c0_n60_w189, 
            w190=> c0_n60_w190, 
            w191=> c0_n60_w191, 
            w192=> c0_n60_w192, 
            w193=> c0_n60_w193, 
            w194=> c0_n60_w194, 
            w195=> c0_n60_w195, 
            w196=> c0_n60_w196, 
            w197=> c0_n60_w197, 
            w198=> c0_n60_w198, 
            w199=> c0_n60_w199, 
            w200=> c0_n60_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n60_y
   );           
            
neuron_inst_61: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n61_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n61_w1, 
            w2=> c0_n61_w2, 
            w3=> c0_n61_w3, 
            w4=> c0_n61_w4, 
            w5=> c0_n61_w5, 
            w6=> c0_n61_w6, 
            w7=> c0_n61_w7, 
            w8=> c0_n61_w8, 
            w9=> c0_n61_w9, 
            w10=> c0_n61_w10, 
            w11=> c0_n61_w11, 
            w12=> c0_n61_w12, 
            w13=> c0_n61_w13, 
            w14=> c0_n61_w14, 
            w15=> c0_n61_w15, 
            w16=> c0_n61_w16, 
            w17=> c0_n61_w17, 
            w18=> c0_n61_w18, 
            w19=> c0_n61_w19, 
            w20=> c0_n61_w20, 
            w21=> c0_n61_w21, 
            w22=> c0_n61_w22, 
            w23=> c0_n61_w23, 
            w24=> c0_n61_w24, 
            w25=> c0_n61_w25, 
            w26=> c0_n61_w26, 
            w27=> c0_n61_w27, 
            w28=> c0_n61_w28, 
            w29=> c0_n61_w29, 
            w30=> c0_n61_w30, 
            w31=> c0_n61_w31, 
            w32=> c0_n61_w32, 
            w33=> c0_n61_w33, 
            w34=> c0_n61_w34, 
            w35=> c0_n61_w35, 
            w36=> c0_n61_w36, 
            w37=> c0_n61_w37, 
            w38=> c0_n61_w38, 
            w39=> c0_n61_w39, 
            w40=> c0_n61_w40, 
            w41=> c0_n61_w41, 
            w42=> c0_n61_w42, 
            w43=> c0_n61_w43, 
            w44=> c0_n61_w44, 
            w45=> c0_n61_w45, 
            w46=> c0_n61_w46, 
            w47=> c0_n61_w47, 
            w48=> c0_n61_w48, 
            w49=> c0_n61_w49, 
            w50=> c0_n61_w50, 
            w51=> c0_n61_w51, 
            w52=> c0_n61_w52, 
            w53=> c0_n61_w53, 
            w54=> c0_n61_w54, 
            w55=> c0_n61_w55, 
            w56=> c0_n61_w56, 
            w57=> c0_n61_w57, 
            w58=> c0_n61_w58, 
            w59=> c0_n61_w59, 
            w60=> c0_n61_w60, 
            w61=> c0_n61_w61, 
            w62=> c0_n61_w62, 
            w63=> c0_n61_w63, 
            w64=> c0_n61_w64, 
            w65=> c0_n61_w65, 
            w66=> c0_n61_w66, 
            w67=> c0_n61_w67, 
            w68=> c0_n61_w68, 
            w69=> c0_n61_w69, 
            w70=> c0_n61_w70, 
            w71=> c0_n61_w71, 
            w72=> c0_n61_w72, 
            w73=> c0_n61_w73, 
            w74=> c0_n61_w74, 
            w75=> c0_n61_w75, 
            w76=> c0_n61_w76, 
            w77=> c0_n61_w77, 
            w78=> c0_n61_w78, 
            w79=> c0_n61_w79, 
            w80=> c0_n61_w80, 
            w81=> c0_n61_w81, 
            w82=> c0_n61_w82, 
            w83=> c0_n61_w83, 
            w84=> c0_n61_w84, 
            w85=> c0_n61_w85, 
            w86=> c0_n61_w86, 
            w87=> c0_n61_w87, 
            w88=> c0_n61_w88, 
            w89=> c0_n61_w89, 
            w90=> c0_n61_w90, 
            w91=> c0_n61_w91, 
            w92=> c0_n61_w92, 
            w93=> c0_n61_w93, 
            w94=> c0_n61_w94, 
            w95=> c0_n61_w95, 
            w96=> c0_n61_w96, 
            w97=> c0_n61_w97, 
            w98=> c0_n61_w98, 
            w99=> c0_n61_w99, 
            w100=> c0_n61_w100, 
            w101=> c0_n61_w101, 
            w102=> c0_n61_w102, 
            w103=> c0_n61_w103, 
            w104=> c0_n61_w104, 
            w105=> c0_n61_w105, 
            w106=> c0_n61_w106, 
            w107=> c0_n61_w107, 
            w108=> c0_n61_w108, 
            w109=> c0_n61_w109, 
            w110=> c0_n61_w110, 
            w111=> c0_n61_w111, 
            w112=> c0_n61_w112, 
            w113=> c0_n61_w113, 
            w114=> c0_n61_w114, 
            w115=> c0_n61_w115, 
            w116=> c0_n61_w116, 
            w117=> c0_n61_w117, 
            w118=> c0_n61_w118, 
            w119=> c0_n61_w119, 
            w120=> c0_n61_w120, 
            w121=> c0_n61_w121, 
            w122=> c0_n61_w122, 
            w123=> c0_n61_w123, 
            w124=> c0_n61_w124, 
            w125=> c0_n61_w125, 
            w126=> c0_n61_w126, 
            w127=> c0_n61_w127, 
            w128=> c0_n61_w128, 
            w129=> c0_n61_w129, 
            w130=> c0_n61_w130, 
            w131=> c0_n61_w131, 
            w132=> c0_n61_w132, 
            w133=> c0_n61_w133, 
            w134=> c0_n61_w134, 
            w135=> c0_n61_w135, 
            w136=> c0_n61_w136, 
            w137=> c0_n61_w137, 
            w138=> c0_n61_w138, 
            w139=> c0_n61_w139, 
            w140=> c0_n61_w140, 
            w141=> c0_n61_w141, 
            w142=> c0_n61_w142, 
            w143=> c0_n61_w143, 
            w144=> c0_n61_w144, 
            w145=> c0_n61_w145, 
            w146=> c0_n61_w146, 
            w147=> c0_n61_w147, 
            w148=> c0_n61_w148, 
            w149=> c0_n61_w149, 
            w150=> c0_n61_w150, 
            w151=> c0_n61_w151, 
            w152=> c0_n61_w152, 
            w153=> c0_n61_w153, 
            w154=> c0_n61_w154, 
            w155=> c0_n61_w155, 
            w156=> c0_n61_w156, 
            w157=> c0_n61_w157, 
            w158=> c0_n61_w158, 
            w159=> c0_n61_w159, 
            w160=> c0_n61_w160, 
            w161=> c0_n61_w161, 
            w162=> c0_n61_w162, 
            w163=> c0_n61_w163, 
            w164=> c0_n61_w164, 
            w165=> c0_n61_w165, 
            w166=> c0_n61_w166, 
            w167=> c0_n61_w167, 
            w168=> c0_n61_w168, 
            w169=> c0_n61_w169, 
            w170=> c0_n61_w170, 
            w171=> c0_n61_w171, 
            w172=> c0_n61_w172, 
            w173=> c0_n61_w173, 
            w174=> c0_n61_w174, 
            w175=> c0_n61_w175, 
            w176=> c0_n61_w176, 
            w177=> c0_n61_w177, 
            w178=> c0_n61_w178, 
            w179=> c0_n61_w179, 
            w180=> c0_n61_w180, 
            w181=> c0_n61_w181, 
            w182=> c0_n61_w182, 
            w183=> c0_n61_w183, 
            w184=> c0_n61_w184, 
            w185=> c0_n61_w185, 
            w186=> c0_n61_w186, 
            w187=> c0_n61_w187, 
            w188=> c0_n61_w188, 
            w189=> c0_n61_w189, 
            w190=> c0_n61_w190, 
            w191=> c0_n61_w191, 
            w192=> c0_n61_w192, 
            w193=> c0_n61_w193, 
            w194=> c0_n61_w194, 
            w195=> c0_n61_w195, 
            w196=> c0_n61_w196, 
            w197=> c0_n61_w197, 
            w198=> c0_n61_w198, 
            w199=> c0_n61_w199, 
            w200=> c0_n61_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n61_y
   );           
            
neuron_inst_62: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n62_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n62_w1, 
            w2=> c0_n62_w2, 
            w3=> c0_n62_w3, 
            w4=> c0_n62_w4, 
            w5=> c0_n62_w5, 
            w6=> c0_n62_w6, 
            w7=> c0_n62_w7, 
            w8=> c0_n62_w8, 
            w9=> c0_n62_w9, 
            w10=> c0_n62_w10, 
            w11=> c0_n62_w11, 
            w12=> c0_n62_w12, 
            w13=> c0_n62_w13, 
            w14=> c0_n62_w14, 
            w15=> c0_n62_w15, 
            w16=> c0_n62_w16, 
            w17=> c0_n62_w17, 
            w18=> c0_n62_w18, 
            w19=> c0_n62_w19, 
            w20=> c0_n62_w20, 
            w21=> c0_n62_w21, 
            w22=> c0_n62_w22, 
            w23=> c0_n62_w23, 
            w24=> c0_n62_w24, 
            w25=> c0_n62_w25, 
            w26=> c0_n62_w26, 
            w27=> c0_n62_w27, 
            w28=> c0_n62_w28, 
            w29=> c0_n62_w29, 
            w30=> c0_n62_w30, 
            w31=> c0_n62_w31, 
            w32=> c0_n62_w32, 
            w33=> c0_n62_w33, 
            w34=> c0_n62_w34, 
            w35=> c0_n62_w35, 
            w36=> c0_n62_w36, 
            w37=> c0_n62_w37, 
            w38=> c0_n62_w38, 
            w39=> c0_n62_w39, 
            w40=> c0_n62_w40, 
            w41=> c0_n62_w41, 
            w42=> c0_n62_w42, 
            w43=> c0_n62_w43, 
            w44=> c0_n62_w44, 
            w45=> c0_n62_w45, 
            w46=> c0_n62_w46, 
            w47=> c0_n62_w47, 
            w48=> c0_n62_w48, 
            w49=> c0_n62_w49, 
            w50=> c0_n62_w50, 
            w51=> c0_n62_w51, 
            w52=> c0_n62_w52, 
            w53=> c0_n62_w53, 
            w54=> c0_n62_w54, 
            w55=> c0_n62_w55, 
            w56=> c0_n62_w56, 
            w57=> c0_n62_w57, 
            w58=> c0_n62_w58, 
            w59=> c0_n62_w59, 
            w60=> c0_n62_w60, 
            w61=> c0_n62_w61, 
            w62=> c0_n62_w62, 
            w63=> c0_n62_w63, 
            w64=> c0_n62_w64, 
            w65=> c0_n62_w65, 
            w66=> c0_n62_w66, 
            w67=> c0_n62_w67, 
            w68=> c0_n62_w68, 
            w69=> c0_n62_w69, 
            w70=> c0_n62_w70, 
            w71=> c0_n62_w71, 
            w72=> c0_n62_w72, 
            w73=> c0_n62_w73, 
            w74=> c0_n62_w74, 
            w75=> c0_n62_w75, 
            w76=> c0_n62_w76, 
            w77=> c0_n62_w77, 
            w78=> c0_n62_w78, 
            w79=> c0_n62_w79, 
            w80=> c0_n62_w80, 
            w81=> c0_n62_w81, 
            w82=> c0_n62_w82, 
            w83=> c0_n62_w83, 
            w84=> c0_n62_w84, 
            w85=> c0_n62_w85, 
            w86=> c0_n62_w86, 
            w87=> c0_n62_w87, 
            w88=> c0_n62_w88, 
            w89=> c0_n62_w89, 
            w90=> c0_n62_w90, 
            w91=> c0_n62_w91, 
            w92=> c0_n62_w92, 
            w93=> c0_n62_w93, 
            w94=> c0_n62_w94, 
            w95=> c0_n62_w95, 
            w96=> c0_n62_w96, 
            w97=> c0_n62_w97, 
            w98=> c0_n62_w98, 
            w99=> c0_n62_w99, 
            w100=> c0_n62_w100, 
            w101=> c0_n62_w101, 
            w102=> c0_n62_w102, 
            w103=> c0_n62_w103, 
            w104=> c0_n62_w104, 
            w105=> c0_n62_w105, 
            w106=> c0_n62_w106, 
            w107=> c0_n62_w107, 
            w108=> c0_n62_w108, 
            w109=> c0_n62_w109, 
            w110=> c0_n62_w110, 
            w111=> c0_n62_w111, 
            w112=> c0_n62_w112, 
            w113=> c0_n62_w113, 
            w114=> c0_n62_w114, 
            w115=> c0_n62_w115, 
            w116=> c0_n62_w116, 
            w117=> c0_n62_w117, 
            w118=> c0_n62_w118, 
            w119=> c0_n62_w119, 
            w120=> c0_n62_w120, 
            w121=> c0_n62_w121, 
            w122=> c0_n62_w122, 
            w123=> c0_n62_w123, 
            w124=> c0_n62_w124, 
            w125=> c0_n62_w125, 
            w126=> c0_n62_w126, 
            w127=> c0_n62_w127, 
            w128=> c0_n62_w128, 
            w129=> c0_n62_w129, 
            w130=> c0_n62_w130, 
            w131=> c0_n62_w131, 
            w132=> c0_n62_w132, 
            w133=> c0_n62_w133, 
            w134=> c0_n62_w134, 
            w135=> c0_n62_w135, 
            w136=> c0_n62_w136, 
            w137=> c0_n62_w137, 
            w138=> c0_n62_w138, 
            w139=> c0_n62_w139, 
            w140=> c0_n62_w140, 
            w141=> c0_n62_w141, 
            w142=> c0_n62_w142, 
            w143=> c0_n62_w143, 
            w144=> c0_n62_w144, 
            w145=> c0_n62_w145, 
            w146=> c0_n62_w146, 
            w147=> c0_n62_w147, 
            w148=> c0_n62_w148, 
            w149=> c0_n62_w149, 
            w150=> c0_n62_w150, 
            w151=> c0_n62_w151, 
            w152=> c0_n62_w152, 
            w153=> c0_n62_w153, 
            w154=> c0_n62_w154, 
            w155=> c0_n62_w155, 
            w156=> c0_n62_w156, 
            w157=> c0_n62_w157, 
            w158=> c0_n62_w158, 
            w159=> c0_n62_w159, 
            w160=> c0_n62_w160, 
            w161=> c0_n62_w161, 
            w162=> c0_n62_w162, 
            w163=> c0_n62_w163, 
            w164=> c0_n62_w164, 
            w165=> c0_n62_w165, 
            w166=> c0_n62_w166, 
            w167=> c0_n62_w167, 
            w168=> c0_n62_w168, 
            w169=> c0_n62_w169, 
            w170=> c0_n62_w170, 
            w171=> c0_n62_w171, 
            w172=> c0_n62_w172, 
            w173=> c0_n62_w173, 
            w174=> c0_n62_w174, 
            w175=> c0_n62_w175, 
            w176=> c0_n62_w176, 
            w177=> c0_n62_w177, 
            w178=> c0_n62_w178, 
            w179=> c0_n62_w179, 
            w180=> c0_n62_w180, 
            w181=> c0_n62_w181, 
            w182=> c0_n62_w182, 
            w183=> c0_n62_w183, 
            w184=> c0_n62_w184, 
            w185=> c0_n62_w185, 
            w186=> c0_n62_w186, 
            w187=> c0_n62_w187, 
            w188=> c0_n62_w188, 
            w189=> c0_n62_w189, 
            w190=> c0_n62_w190, 
            w191=> c0_n62_w191, 
            w192=> c0_n62_w192, 
            w193=> c0_n62_w193, 
            w194=> c0_n62_w194, 
            w195=> c0_n62_w195, 
            w196=> c0_n62_w196, 
            w197=> c0_n62_w197, 
            w198=> c0_n62_w198, 
            w199=> c0_n62_w199, 
            w200=> c0_n62_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n62_y
   );           
            
neuron_inst_63: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n63_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n63_w1, 
            w2=> c0_n63_w2, 
            w3=> c0_n63_w3, 
            w4=> c0_n63_w4, 
            w5=> c0_n63_w5, 
            w6=> c0_n63_w6, 
            w7=> c0_n63_w7, 
            w8=> c0_n63_w8, 
            w9=> c0_n63_w9, 
            w10=> c0_n63_w10, 
            w11=> c0_n63_w11, 
            w12=> c0_n63_w12, 
            w13=> c0_n63_w13, 
            w14=> c0_n63_w14, 
            w15=> c0_n63_w15, 
            w16=> c0_n63_w16, 
            w17=> c0_n63_w17, 
            w18=> c0_n63_w18, 
            w19=> c0_n63_w19, 
            w20=> c0_n63_w20, 
            w21=> c0_n63_w21, 
            w22=> c0_n63_w22, 
            w23=> c0_n63_w23, 
            w24=> c0_n63_w24, 
            w25=> c0_n63_w25, 
            w26=> c0_n63_w26, 
            w27=> c0_n63_w27, 
            w28=> c0_n63_w28, 
            w29=> c0_n63_w29, 
            w30=> c0_n63_w30, 
            w31=> c0_n63_w31, 
            w32=> c0_n63_w32, 
            w33=> c0_n63_w33, 
            w34=> c0_n63_w34, 
            w35=> c0_n63_w35, 
            w36=> c0_n63_w36, 
            w37=> c0_n63_w37, 
            w38=> c0_n63_w38, 
            w39=> c0_n63_w39, 
            w40=> c0_n63_w40, 
            w41=> c0_n63_w41, 
            w42=> c0_n63_w42, 
            w43=> c0_n63_w43, 
            w44=> c0_n63_w44, 
            w45=> c0_n63_w45, 
            w46=> c0_n63_w46, 
            w47=> c0_n63_w47, 
            w48=> c0_n63_w48, 
            w49=> c0_n63_w49, 
            w50=> c0_n63_w50, 
            w51=> c0_n63_w51, 
            w52=> c0_n63_w52, 
            w53=> c0_n63_w53, 
            w54=> c0_n63_w54, 
            w55=> c0_n63_w55, 
            w56=> c0_n63_w56, 
            w57=> c0_n63_w57, 
            w58=> c0_n63_w58, 
            w59=> c0_n63_w59, 
            w60=> c0_n63_w60, 
            w61=> c0_n63_w61, 
            w62=> c0_n63_w62, 
            w63=> c0_n63_w63, 
            w64=> c0_n63_w64, 
            w65=> c0_n63_w65, 
            w66=> c0_n63_w66, 
            w67=> c0_n63_w67, 
            w68=> c0_n63_w68, 
            w69=> c0_n63_w69, 
            w70=> c0_n63_w70, 
            w71=> c0_n63_w71, 
            w72=> c0_n63_w72, 
            w73=> c0_n63_w73, 
            w74=> c0_n63_w74, 
            w75=> c0_n63_w75, 
            w76=> c0_n63_w76, 
            w77=> c0_n63_w77, 
            w78=> c0_n63_w78, 
            w79=> c0_n63_w79, 
            w80=> c0_n63_w80, 
            w81=> c0_n63_w81, 
            w82=> c0_n63_w82, 
            w83=> c0_n63_w83, 
            w84=> c0_n63_w84, 
            w85=> c0_n63_w85, 
            w86=> c0_n63_w86, 
            w87=> c0_n63_w87, 
            w88=> c0_n63_w88, 
            w89=> c0_n63_w89, 
            w90=> c0_n63_w90, 
            w91=> c0_n63_w91, 
            w92=> c0_n63_w92, 
            w93=> c0_n63_w93, 
            w94=> c0_n63_w94, 
            w95=> c0_n63_w95, 
            w96=> c0_n63_w96, 
            w97=> c0_n63_w97, 
            w98=> c0_n63_w98, 
            w99=> c0_n63_w99, 
            w100=> c0_n63_w100, 
            w101=> c0_n63_w101, 
            w102=> c0_n63_w102, 
            w103=> c0_n63_w103, 
            w104=> c0_n63_w104, 
            w105=> c0_n63_w105, 
            w106=> c0_n63_w106, 
            w107=> c0_n63_w107, 
            w108=> c0_n63_w108, 
            w109=> c0_n63_w109, 
            w110=> c0_n63_w110, 
            w111=> c0_n63_w111, 
            w112=> c0_n63_w112, 
            w113=> c0_n63_w113, 
            w114=> c0_n63_w114, 
            w115=> c0_n63_w115, 
            w116=> c0_n63_w116, 
            w117=> c0_n63_w117, 
            w118=> c0_n63_w118, 
            w119=> c0_n63_w119, 
            w120=> c0_n63_w120, 
            w121=> c0_n63_w121, 
            w122=> c0_n63_w122, 
            w123=> c0_n63_w123, 
            w124=> c0_n63_w124, 
            w125=> c0_n63_w125, 
            w126=> c0_n63_w126, 
            w127=> c0_n63_w127, 
            w128=> c0_n63_w128, 
            w129=> c0_n63_w129, 
            w130=> c0_n63_w130, 
            w131=> c0_n63_w131, 
            w132=> c0_n63_w132, 
            w133=> c0_n63_w133, 
            w134=> c0_n63_w134, 
            w135=> c0_n63_w135, 
            w136=> c0_n63_w136, 
            w137=> c0_n63_w137, 
            w138=> c0_n63_w138, 
            w139=> c0_n63_w139, 
            w140=> c0_n63_w140, 
            w141=> c0_n63_w141, 
            w142=> c0_n63_w142, 
            w143=> c0_n63_w143, 
            w144=> c0_n63_w144, 
            w145=> c0_n63_w145, 
            w146=> c0_n63_w146, 
            w147=> c0_n63_w147, 
            w148=> c0_n63_w148, 
            w149=> c0_n63_w149, 
            w150=> c0_n63_w150, 
            w151=> c0_n63_w151, 
            w152=> c0_n63_w152, 
            w153=> c0_n63_w153, 
            w154=> c0_n63_w154, 
            w155=> c0_n63_w155, 
            w156=> c0_n63_w156, 
            w157=> c0_n63_w157, 
            w158=> c0_n63_w158, 
            w159=> c0_n63_w159, 
            w160=> c0_n63_w160, 
            w161=> c0_n63_w161, 
            w162=> c0_n63_w162, 
            w163=> c0_n63_w163, 
            w164=> c0_n63_w164, 
            w165=> c0_n63_w165, 
            w166=> c0_n63_w166, 
            w167=> c0_n63_w167, 
            w168=> c0_n63_w168, 
            w169=> c0_n63_w169, 
            w170=> c0_n63_w170, 
            w171=> c0_n63_w171, 
            w172=> c0_n63_w172, 
            w173=> c0_n63_w173, 
            w174=> c0_n63_w174, 
            w175=> c0_n63_w175, 
            w176=> c0_n63_w176, 
            w177=> c0_n63_w177, 
            w178=> c0_n63_w178, 
            w179=> c0_n63_w179, 
            w180=> c0_n63_w180, 
            w181=> c0_n63_w181, 
            w182=> c0_n63_w182, 
            w183=> c0_n63_w183, 
            w184=> c0_n63_w184, 
            w185=> c0_n63_w185, 
            w186=> c0_n63_w186, 
            w187=> c0_n63_w187, 
            w188=> c0_n63_w188, 
            w189=> c0_n63_w189, 
            w190=> c0_n63_w190, 
            w191=> c0_n63_w191, 
            w192=> c0_n63_w192, 
            w193=> c0_n63_w193, 
            w194=> c0_n63_w194, 
            w195=> c0_n63_w195, 
            w196=> c0_n63_w196, 
            w197=> c0_n63_w197, 
            w198=> c0_n63_w198, 
            w199=> c0_n63_w199, 
            w200=> c0_n63_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n63_y
   );           
            
neuron_inst_64: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n64_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n64_w1, 
            w2=> c0_n64_w2, 
            w3=> c0_n64_w3, 
            w4=> c0_n64_w4, 
            w5=> c0_n64_w5, 
            w6=> c0_n64_w6, 
            w7=> c0_n64_w7, 
            w8=> c0_n64_w8, 
            w9=> c0_n64_w9, 
            w10=> c0_n64_w10, 
            w11=> c0_n64_w11, 
            w12=> c0_n64_w12, 
            w13=> c0_n64_w13, 
            w14=> c0_n64_w14, 
            w15=> c0_n64_w15, 
            w16=> c0_n64_w16, 
            w17=> c0_n64_w17, 
            w18=> c0_n64_w18, 
            w19=> c0_n64_w19, 
            w20=> c0_n64_w20, 
            w21=> c0_n64_w21, 
            w22=> c0_n64_w22, 
            w23=> c0_n64_w23, 
            w24=> c0_n64_w24, 
            w25=> c0_n64_w25, 
            w26=> c0_n64_w26, 
            w27=> c0_n64_w27, 
            w28=> c0_n64_w28, 
            w29=> c0_n64_w29, 
            w30=> c0_n64_w30, 
            w31=> c0_n64_w31, 
            w32=> c0_n64_w32, 
            w33=> c0_n64_w33, 
            w34=> c0_n64_w34, 
            w35=> c0_n64_w35, 
            w36=> c0_n64_w36, 
            w37=> c0_n64_w37, 
            w38=> c0_n64_w38, 
            w39=> c0_n64_w39, 
            w40=> c0_n64_w40, 
            w41=> c0_n64_w41, 
            w42=> c0_n64_w42, 
            w43=> c0_n64_w43, 
            w44=> c0_n64_w44, 
            w45=> c0_n64_w45, 
            w46=> c0_n64_w46, 
            w47=> c0_n64_w47, 
            w48=> c0_n64_w48, 
            w49=> c0_n64_w49, 
            w50=> c0_n64_w50, 
            w51=> c0_n64_w51, 
            w52=> c0_n64_w52, 
            w53=> c0_n64_w53, 
            w54=> c0_n64_w54, 
            w55=> c0_n64_w55, 
            w56=> c0_n64_w56, 
            w57=> c0_n64_w57, 
            w58=> c0_n64_w58, 
            w59=> c0_n64_w59, 
            w60=> c0_n64_w60, 
            w61=> c0_n64_w61, 
            w62=> c0_n64_w62, 
            w63=> c0_n64_w63, 
            w64=> c0_n64_w64, 
            w65=> c0_n64_w65, 
            w66=> c0_n64_w66, 
            w67=> c0_n64_w67, 
            w68=> c0_n64_w68, 
            w69=> c0_n64_w69, 
            w70=> c0_n64_w70, 
            w71=> c0_n64_w71, 
            w72=> c0_n64_w72, 
            w73=> c0_n64_w73, 
            w74=> c0_n64_w74, 
            w75=> c0_n64_w75, 
            w76=> c0_n64_w76, 
            w77=> c0_n64_w77, 
            w78=> c0_n64_w78, 
            w79=> c0_n64_w79, 
            w80=> c0_n64_w80, 
            w81=> c0_n64_w81, 
            w82=> c0_n64_w82, 
            w83=> c0_n64_w83, 
            w84=> c0_n64_w84, 
            w85=> c0_n64_w85, 
            w86=> c0_n64_w86, 
            w87=> c0_n64_w87, 
            w88=> c0_n64_w88, 
            w89=> c0_n64_w89, 
            w90=> c0_n64_w90, 
            w91=> c0_n64_w91, 
            w92=> c0_n64_w92, 
            w93=> c0_n64_w93, 
            w94=> c0_n64_w94, 
            w95=> c0_n64_w95, 
            w96=> c0_n64_w96, 
            w97=> c0_n64_w97, 
            w98=> c0_n64_w98, 
            w99=> c0_n64_w99, 
            w100=> c0_n64_w100, 
            w101=> c0_n64_w101, 
            w102=> c0_n64_w102, 
            w103=> c0_n64_w103, 
            w104=> c0_n64_w104, 
            w105=> c0_n64_w105, 
            w106=> c0_n64_w106, 
            w107=> c0_n64_w107, 
            w108=> c0_n64_w108, 
            w109=> c0_n64_w109, 
            w110=> c0_n64_w110, 
            w111=> c0_n64_w111, 
            w112=> c0_n64_w112, 
            w113=> c0_n64_w113, 
            w114=> c0_n64_w114, 
            w115=> c0_n64_w115, 
            w116=> c0_n64_w116, 
            w117=> c0_n64_w117, 
            w118=> c0_n64_w118, 
            w119=> c0_n64_w119, 
            w120=> c0_n64_w120, 
            w121=> c0_n64_w121, 
            w122=> c0_n64_w122, 
            w123=> c0_n64_w123, 
            w124=> c0_n64_w124, 
            w125=> c0_n64_w125, 
            w126=> c0_n64_w126, 
            w127=> c0_n64_w127, 
            w128=> c0_n64_w128, 
            w129=> c0_n64_w129, 
            w130=> c0_n64_w130, 
            w131=> c0_n64_w131, 
            w132=> c0_n64_w132, 
            w133=> c0_n64_w133, 
            w134=> c0_n64_w134, 
            w135=> c0_n64_w135, 
            w136=> c0_n64_w136, 
            w137=> c0_n64_w137, 
            w138=> c0_n64_w138, 
            w139=> c0_n64_w139, 
            w140=> c0_n64_w140, 
            w141=> c0_n64_w141, 
            w142=> c0_n64_w142, 
            w143=> c0_n64_w143, 
            w144=> c0_n64_w144, 
            w145=> c0_n64_w145, 
            w146=> c0_n64_w146, 
            w147=> c0_n64_w147, 
            w148=> c0_n64_w148, 
            w149=> c0_n64_w149, 
            w150=> c0_n64_w150, 
            w151=> c0_n64_w151, 
            w152=> c0_n64_w152, 
            w153=> c0_n64_w153, 
            w154=> c0_n64_w154, 
            w155=> c0_n64_w155, 
            w156=> c0_n64_w156, 
            w157=> c0_n64_w157, 
            w158=> c0_n64_w158, 
            w159=> c0_n64_w159, 
            w160=> c0_n64_w160, 
            w161=> c0_n64_w161, 
            w162=> c0_n64_w162, 
            w163=> c0_n64_w163, 
            w164=> c0_n64_w164, 
            w165=> c0_n64_w165, 
            w166=> c0_n64_w166, 
            w167=> c0_n64_w167, 
            w168=> c0_n64_w168, 
            w169=> c0_n64_w169, 
            w170=> c0_n64_w170, 
            w171=> c0_n64_w171, 
            w172=> c0_n64_w172, 
            w173=> c0_n64_w173, 
            w174=> c0_n64_w174, 
            w175=> c0_n64_w175, 
            w176=> c0_n64_w176, 
            w177=> c0_n64_w177, 
            w178=> c0_n64_w178, 
            w179=> c0_n64_w179, 
            w180=> c0_n64_w180, 
            w181=> c0_n64_w181, 
            w182=> c0_n64_w182, 
            w183=> c0_n64_w183, 
            w184=> c0_n64_w184, 
            w185=> c0_n64_w185, 
            w186=> c0_n64_w186, 
            w187=> c0_n64_w187, 
            w188=> c0_n64_w188, 
            w189=> c0_n64_w189, 
            w190=> c0_n64_w190, 
            w191=> c0_n64_w191, 
            w192=> c0_n64_w192, 
            w193=> c0_n64_w193, 
            w194=> c0_n64_w194, 
            w195=> c0_n64_w195, 
            w196=> c0_n64_w196, 
            w197=> c0_n64_w197, 
            w198=> c0_n64_w198, 
            w199=> c0_n64_w199, 
            w200=> c0_n64_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n64_y
   );           
            
neuron_inst_65: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n65_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n65_w1, 
            w2=> c0_n65_w2, 
            w3=> c0_n65_w3, 
            w4=> c0_n65_w4, 
            w5=> c0_n65_w5, 
            w6=> c0_n65_w6, 
            w7=> c0_n65_w7, 
            w8=> c0_n65_w8, 
            w9=> c0_n65_w9, 
            w10=> c0_n65_w10, 
            w11=> c0_n65_w11, 
            w12=> c0_n65_w12, 
            w13=> c0_n65_w13, 
            w14=> c0_n65_w14, 
            w15=> c0_n65_w15, 
            w16=> c0_n65_w16, 
            w17=> c0_n65_w17, 
            w18=> c0_n65_w18, 
            w19=> c0_n65_w19, 
            w20=> c0_n65_w20, 
            w21=> c0_n65_w21, 
            w22=> c0_n65_w22, 
            w23=> c0_n65_w23, 
            w24=> c0_n65_w24, 
            w25=> c0_n65_w25, 
            w26=> c0_n65_w26, 
            w27=> c0_n65_w27, 
            w28=> c0_n65_w28, 
            w29=> c0_n65_w29, 
            w30=> c0_n65_w30, 
            w31=> c0_n65_w31, 
            w32=> c0_n65_w32, 
            w33=> c0_n65_w33, 
            w34=> c0_n65_w34, 
            w35=> c0_n65_w35, 
            w36=> c0_n65_w36, 
            w37=> c0_n65_w37, 
            w38=> c0_n65_w38, 
            w39=> c0_n65_w39, 
            w40=> c0_n65_w40, 
            w41=> c0_n65_w41, 
            w42=> c0_n65_w42, 
            w43=> c0_n65_w43, 
            w44=> c0_n65_w44, 
            w45=> c0_n65_w45, 
            w46=> c0_n65_w46, 
            w47=> c0_n65_w47, 
            w48=> c0_n65_w48, 
            w49=> c0_n65_w49, 
            w50=> c0_n65_w50, 
            w51=> c0_n65_w51, 
            w52=> c0_n65_w52, 
            w53=> c0_n65_w53, 
            w54=> c0_n65_w54, 
            w55=> c0_n65_w55, 
            w56=> c0_n65_w56, 
            w57=> c0_n65_w57, 
            w58=> c0_n65_w58, 
            w59=> c0_n65_w59, 
            w60=> c0_n65_w60, 
            w61=> c0_n65_w61, 
            w62=> c0_n65_w62, 
            w63=> c0_n65_w63, 
            w64=> c0_n65_w64, 
            w65=> c0_n65_w65, 
            w66=> c0_n65_w66, 
            w67=> c0_n65_w67, 
            w68=> c0_n65_w68, 
            w69=> c0_n65_w69, 
            w70=> c0_n65_w70, 
            w71=> c0_n65_w71, 
            w72=> c0_n65_w72, 
            w73=> c0_n65_w73, 
            w74=> c0_n65_w74, 
            w75=> c0_n65_w75, 
            w76=> c0_n65_w76, 
            w77=> c0_n65_w77, 
            w78=> c0_n65_w78, 
            w79=> c0_n65_w79, 
            w80=> c0_n65_w80, 
            w81=> c0_n65_w81, 
            w82=> c0_n65_w82, 
            w83=> c0_n65_w83, 
            w84=> c0_n65_w84, 
            w85=> c0_n65_w85, 
            w86=> c0_n65_w86, 
            w87=> c0_n65_w87, 
            w88=> c0_n65_w88, 
            w89=> c0_n65_w89, 
            w90=> c0_n65_w90, 
            w91=> c0_n65_w91, 
            w92=> c0_n65_w92, 
            w93=> c0_n65_w93, 
            w94=> c0_n65_w94, 
            w95=> c0_n65_w95, 
            w96=> c0_n65_w96, 
            w97=> c0_n65_w97, 
            w98=> c0_n65_w98, 
            w99=> c0_n65_w99, 
            w100=> c0_n65_w100, 
            w101=> c0_n65_w101, 
            w102=> c0_n65_w102, 
            w103=> c0_n65_w103, 
            w104=> c0_n65_w104, 
            w105=> c0_n65_w105, 
            w106=> c0_n65_w106, 
            w107=> c0_n65_w107, 
            w108=> c0_n65_w108, 
            w109=> c0_n65_w109, 
            w110=> c0_n65_w110, 
            w111=> c0_n65_w111, 
            w112=> c0_n65_w112, 
            w113=> c0_n65_w113, 
            w114=> c0_n65_w114, 
            w115=> c0_n65_w115, 
            w116=> c0_n65_w116, 
            w117=> c0_n65_w117, 
            w118=> c0_n65_w118, 
            w119=> c0_n65_w119, 
            w120=> c0_n65_w120, 
            w121=> c0_n65_w121, 
            w122=> c0_n65_w122, 
            w123=> c0_n65_w123, 
            w124=> c0_n65_w124, 
            w125=> c0_n65_w125, 
            w126=> c0_n65_w126, 
            w127=> c0_n65_w127, 
            w128=> c0_n65_w128, 
            w129=> c0_n65_w129, 
            w130=> c0_n65_w130, 
            w131=> c0_n65_w131, 
            w132=> c0_n65_w132, 
            w133=> c0_n65_w133, 
            w134=> c0_n65_w134, 
            w135=> c0_n65_w135, 
            w136=> c0_n65_w136, 
            w137=> c0_n65_w137, 
            w138=> c0_n65_w138, 
            w139=> c0_n65_w139, 
            w140=> c0_n65_w140, 
            w141=> c0_n65_w141, 
            w142=> c0_n65_w142, 
            w143=> c0_n65_w143, 
            w144=> c0_n65_w144, 
            w145=> c0_n65_w145, 
            w146=> c0_n65_w146, 
            w147=> c0_n65_w147, 
            w148=> c0_n65_w148, 
            w149=> c0_n65_w149, 
            w150=> c0_n65_w150, 
            w151=> c0_n65_w151, 
            w152=> c0_n65_w152, 
            w153=> c0_n65_w153, 
            w154=> c0_n65_w154, 
            w155=> c0_n65_w155, 
            w156=> c0_n65_w156, 
            w157=> c0_n65_w157, 
            w158=> c0_n65_w158, 
            w159=> c0_n65_w159, 
            w160=> c0_n65_w160, 
            w161=> c0_n65_w161, 
            w162=> c0_n65_w162, 
            w163=> c0_n65_w163, 
            w164=> c0_n65_w164, 
            w165=> c0_n65_w165, 
            w166=> c0_n65_w166, 
            w167=> c0_n65_w167, 
            w168=> c0_n65_w168, 
            w169=> c0_n65_w169, 
            w170=> c0_n65_w170, 
            w171=> c0_n65_w171, 
            w172=> c0_n65_w172, 
            w173=> c0_n65_w173, 
            w174=> c0_n65_w174, 
            w175=> c0_n65_w175, 
            w176=> c0_n65_w176, 
            w177=> c0_n65_w177, 
            w178=> c0_n65_w178, 
            w179=> c0_n65_w179, 
            w180=> c0_n65_w180, 
            w181=> c0_n65_w181, 
            w182=> c0_n65_w182, 
            w183=> c0_n65_w183, 
            w184=> c0_n65_w184, 
            w185=> c0_n65_w185, 
            w186=> c0_n65_w186, 
            w187=> c0_n65_w187, 
            w188=> c0_n65_w188, 
            w189=> c0_n65_w189, 
            w190=> c0_n65_w190, 
            w191=> c0_n65_w191, 
            w192=> c0_n65_w192, 
            w193=> c0_n65_w193, 
            w194=> c0_n65_w194, 
            w195=> c0_n65_w195, 
            w196=> c0_n65_w196, 
            w197=> c0_n65_w197, 
            w198=> c0_n65_w198, 
            w199=> c0_n65_w199, 
            w200=> c0_n65_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n65_y
   );           
            
neuron_inst_66: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n66_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n66_w1, 
            w2=> c0_n66_w2, 
            w3=> c0_n66_w3, 
            w4=> c0_n66_w4, 
            w5=> c0_n66_w5, 
            w6=> c0_n66_w6, 
            w7=> c0_n66_w7, 
            w8=> c0_n66_w8, 
            w9=> c0_n66_w9, 
            w10=> c0_n66_w10, 
            w11=> c0_n66_w11, 
            w12=> c0_n66_w12, 
            w13=> c0_n66_w13, 
            w14=> c0_n66_w14, 
            w15=> c0_n66_w15, 
            w16=> c0_n66_w16, 
            w17=> c0_n66_w17, 
            w18=> c0_n66_w18, 
            w19=> c0_n66_w19, 
            w20=> c0_n66_w20, 
            w21=> c0_n66_w21, 
            w22=> c0_n66_w22, 
            w23=> c0_n66_w23, 
            w24=> c0_n66_w24, 
            w25=> c0_n66_w25, 
            w26=> c0_n66_w26, 
            w27=> c0_n66_w27, 
            w28=> c0_n66_w28, 
            w29=> c0_n66_w29, 
            w30=> c0_n66_w30, 
            w31=> c0_n66_w31, 
            w32=> c0_n66_w32, 
            w33=> c0_n66_w33, 
            w34=> c0_n66_w34, 
            w35=> c0_n66_w35, 
            w36=> c0_n66_w36, 
            w37=> c0_n66_w37, 
            w38=> c0_n66_w38, 
            w39=> c0_n66_w39, 
            w40=> c0_n66_w40, 
            w41=> c0_n66_w41, 
            w42=> c0_n66_w42, 
            w43=> c0_n66_w43, 
            w44=> c0_n66_w44, 
            w45=> c0_n66_w45, 
            w46=> c0_n66_w46, 
            w47=> c0_n66_w47, 
            w48=> c0_n66_w48, 
            w49=> c0_n66_w49, 
            w50=> c0_n66_w50, 
            w51=> c0_n66_w51, 
            w52=> c0_n66_w52, 
            w53=> c0_n66_w53, 
            w54=> c0_n66_w54, 
            w55=> c0_n66_w55, 
            w56=> c0_n66_w56, 
            w57=> c0_n66_w57, 
            w58=> c0_n66_w58, 
            w59=> c0_n66_w59, 
            w60=> c0_n66_w60, 
            w61=> c0_n66_w61, 
            w62=> c0_n66_w62, 
            w63=> c0_n66_w63, 
            w64=> c0_n66_w64, 
            w65=> c0_n66_w65, 
            w66=> c0_n66_w66, 
            w67=> c0_n66_w67, 
            w68=> c0_n66_w68, 
            w69=> c0_n66_w69, 
            w70=> c0_n66_w70, 
            w71=> c0_n66_w71, 
            w72=> c0_n66_w72, 
            w73=> c0_n66_w73, 
            w74=> c0_n66_w74, 
            w75=> c0_n66_w75, 
            w76=> c0_n66_w76, 
            w77=> c0_n66_w77, 
            w78=> c0_n66_w78, 
            w79=> c0_n66_w79, 
            w80=> c0_n66_w80, 
            w81=> c0_n66_w81, 
            w82=> c0_n66_w82, 
            w83=> c0_n66_w83, 
            w84=> c0_n66_w84, 
            w85=> c0_n66_w85, 
            w86=> c0_n66_w86, 
            w87=> c0_n66_w87, 
            w88=> c0_n66_w88, 
            w89=> c0_n66_w89, 
            w90=> c0_n66_w90, 
            w91=> c0_n66_w91, 
            w92=> c0_n66_w92, 
            w93=> c0_n66_w93, 
            w94=> c0_n66_w94, 
            w95=> c0_n66_w95, 
            w96=> c0_n66_w96, 
            w97=> c0_n66_w97, 
            w98=> c0_n66_w98, 
            w99=> c0_n66_w99, 
            w100=> c0_n66_w100, 
            w101=> c0_n66_w101, 
            w102=> c0_n66_w102, 
            w103=> c0_n66_w103, 
            w104=> c0_n66_w104, 
            w105=> c0_n66_w105, 
            w106=> c0_n66_w106, 
            w107=> c0_n66_w107, 
            w108=> c0_n66_w108, 
            w109=> c0_n66_w109, 
            w110=> c0_n66_w110, 
            w111=> c0_n66_w111, 
            w112=> c0_n66_w112, 
            w113=> c0_n66_w113, 
            w114=> c0_n66_w114, 
            w115=> c0_n66_w115, 
            w116=> c0_n66_w116, 
            w117=> c0_n66_w117, 
            w118=> c0_n66_w118, 
            w119=> c0_n66_w119, 
            w120=> c0_n66_w120, 
            w121=> c0_n66_w121, 
            w122=> c0_n66_w122, 
            w123=> c0_n66_w123, 
            w124=> c0_n66_w124, 
            w125=> c0_n66_w125, 
            w126=> c0_n66_w126, 
            w127=> c0_n66_w127, 
            w128=> c0_n66_w128, 
            w129=> c0_n66_w129, 
            w130=> c0_n66_w130, 
            w131=> c0_n66_w131, 
            w132=> c0_n66_w132, 
            w133=> c0_n66_w133, 
            w134=> c0_n66_w134, 
            w135=> c0_n66_w135, 
            w136=> c0_n66_w136, 
            w137=> c0_n66_w137, 
            w138=> c0_n66_w138, 
            w139=> c0_n66_w139, 
            w140=> c0_n66_w140, 
            w141=> c0_n66_w141, 
            w142=> c0_n66_w142, 
            w143=> c0_n66_w143, 
            w144=> c0_n66_w144, 
            w145=> c0_n66_w145, 
            w146=> c0_n66_w146, 
            w147=> c0_n66_w147, 
            w148=> c0_n66_w148, 
            w149=> c0_n66_w149, 
            w150=> c0_n66_w150, 
            w151=> c0_n66_w151, 
            w152=> c0_n66_w152, 
            w153=> c0_n66_w153, 
            w154=> c0_n66_w154, 
            w155=> c0_n66_w155, 
            w156=> c0_n66_w156, 
            w157=> c0_n66_w157, 
            w158=> c0_n66_w158, 
            w159=> c0_n66_w159, 
            w160=> c0_n66_w160, 
            w161=> c0_n66_w161, 
            w162=> c0_n66_w162, 
            w163=> c0_n66_w163, 
            w164=> c0_n66_w164, 
            w165=> c0_n66_w165, 
            w166=> c0_n66_w166, 
            w167=> c0_n66_w167, 
            w168=> c0_n66_w168, 
            w169=> c0_n66_w169, 
            w170=> c0_n66_w170, 
            w171=> c0_n66_w171, 
            w172=> c0_n66_w172, 
            w173=> c0_n66_w173, 
            w174=> c0_n66_w174, 
            w175=> c0_n66_w175, 
            w176=> c0_n66_w176, 
            w177=> c0_n66_w177, 
            w178=> c0_n66_w178, 
            w179=> c0_n66_w179, 
            w180=> c0_n66_w180, 
            w181=> c0_n66_w181, 
            w182=> c0_n66_w182, 
            w183=> c0_n66_w183, 
            w184=> c0_n66_w184, 
            w185=> c0_n66_w185, 
            w186=> c0_n66_w186, 
            w187=> c0_n66_w187, 
            w188=> c0_n66_w188, 
            w189=> c0_n66_w189, 
            w190=> c0_n66_w190, 
            w191=> c0_n66_w191, 
            w192=> c0_n66_w192, 
            w193=> c0_n66_w193, 
            w194=> c0_n66_w194, 
            w195=> c0_n66_w195, 
            w196=> c0_n66_w196, 
            w197=> c0_n66_w197, 
            w198=> c0_n66_w198, 
            w199=> c0_n66_w199, 
            w200=> c0_n66_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n66_y
   );           
            
neuron_inst_67: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n67_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n67_w1, 
            w2=> c0_n67_w2, 
            w3=> c0_n67_w3, 
            w4=> c0_n67_w4, 
            w5=> c0_n67_w5, 
            w6=> c0_n67_w6, 
            w7=> c0_n67_w7, 
            w8=> c0_n67_w8, 
            w9=> c0_n67_w9, 
            w10=> c0_n67_w10, 
            w11=> c0_n67_w11, 
            w12=> c0_n67_w12, 
            w13=> c0_n67_w13, 
            w14=> c0_n67_w14, 
            w15=> c0_n67_w15, 
            w16=> c0_n67_w16, 
            w17=> c0_n67_w17, 
            w18=> c0_n67_w18, 
            w19=> c0_n67_w19, 
            w20=> c0_n67_w20, 
            w21=> c0_n67_w21, 
            w22=> c0_n67_w22, 
            w23=> c0_n67_w23, 
            w24=> c0_n67_w24, 
            w25=> c0_n67_w25, 
            w26=> c0_n67_w26, 
            w27=> c0_n67_w27, 
            w28=> c0_n67_w28, 
            w29=> c0_n67_w29, 
            w30=> c0_n67_w30, 
            w31=> c0_n67_w31, 
            w32=> c0_n67_w32, 
            w33=> c0_n67_w33, 
            w34=> c0_n67_w34, 
            w35=> c0_n67_w35, 
            w36=> c0_n67_w36, 
            w37=> c0_n67_w37, 
            w38=> c0_n67_w38, 
            w39=> c0_n67_w39, 
            w40=> c0_n67_w40, 
            w41=> c0_n67_w41, 
            w42=> c0_n67_w42, 
            w43=> c0_n67_w43, 
            w44=> c0_n67_w44, 
            w45=> c0_n67_w45, 
            w46=> c0_n67_w46, 
            w47=> c0_n67_w47, 
            w48=> c0_n67_w48, 
            w49=> c0_n67_w49, 
            w50=> c0_n67_w50, 
            w51=> c0_n67_w51, 
            w52=> c0_n67_w52, 
            w53=> c0_n67_w53, 
            w54=> c0_n67_w54, 
            w55=> c0_n67_w55, 
            w56=> c0_n67_w56, 
            w57=> c0_n67_w57, 
            w58=> c0_n67_w58, 
            w59=> c0_n67_w59, 
            w60=> c0_n67_w60, 
            w61=> c0_n67_w61, 
            w62=> c0_n67_w62, 
            w63=> c0_n67_w63, 
            w64=> c0_n67_w64, 
            w65=> c0_n67_w65, 
            w66=> c0_n67_w66, 
            w67=> c0_n67_w67, 
            w68=> c0_n67_w68, 
            w69=> c0_n67_w69, 
            w70=> c0_n67_w70, 
            w71=> c0_n67_w71, 
            w72=> c0_n67_w72, 
            w73=> c0_n67_w73, 
            w74=> c0_n67_w74, 
            w75=> c0_n67_w75, 
            w76=> c0_n67_w76, 
            w77=> c0_n67_w77, 
            w78=> c0_n67_w78, 
            w79=> c0_n67_w79, 
            w80=> c0_n67_w80, 
            w81=> c0_n67_w81, 
            w82=> c0_n67_w82, 
            w83=> c0_n67_w83, 
            w84=> c0_n67_w84, 
            w85=> c0_n67_w85, 
            w86=> c0_n67_w86, 
            w87=> c0_n67_w87, 
            w88=> c0_n67_w88, 
            w89=> c0_n67_w89, 
            w90=> c0_n67_w90, 
            w91=> c0_n67_w91, 
            w92=> c0_n67_w92, 
            w93=> c0_n67_w93, 
            w94=> c0_n67_w94, 
            w95=> c0_n67_w95, 
            w96=> c0_n67_w96, 
            w97=> c0_n67_w97, 
            w98=> c0_n67_w98, 
            w99=> c0_n67_w99, 
            w100=> c0_n67_w100, 
            w101=> c0_n67_w101, 
            w102=> c0_n67_w102, 
            w103=> c0_n67_w103, 
            w104=> c0_n67_w104, 
            w105=> c0_n67_w105, 
            w106=> c0_n67_w106, 
            w107=> c0_n67_w107, 
            w108=> c0_n67_w108, 
            w109=> c0_n67_w109, 
            w110=> c0_n67_w110, 
            w111=> c0_n67_w111, 
            w112=> c0_n67_w112, 
            w113=> c0_n67_w113, 
            w114=> c0_n67_w114, 
            w115=> c0_n67_w115, 
            w116=> c0_n67_w116, 
            w117=> c0_n67_w117, 
            w118=> c0_n67_w118, 
            w119=> c0_n67_w119, 
            w120=> c0_n67_w120, 
            w121=> c0_n67_w121, 
            w122=> c0_n67_w122, 
            w123=> c0_n67_w123, 
            w124=> c0_n67_w124, 
            w125=> c0_n67_w125, 
            w126=> c0_n67_w126, 
            w127=> c0_n67_w127, 
            w128=> c0_n67_w128, 
            w129=> c0_n67_w129, 
            w130=> c0_n67_w130, 
            w131=> c0_n67_w131, 
            w132=> c0_n67_w132, 
            w133=> c0_n67_w133, 
            w134=> c0_n67_w134, 
            w135=> c0_n67_w135, 
            w136=> c0_n67_w136, 
            w137=> c0_n67_w137, 
            w138=> c0_n67_w138, 
            w139=> c0_n67_w139, 
            w140=> c0_n67_w140, 
            w141=> c0_n67_w141, 
            w142=> c0_n67_w142, 
            w143=> c0_n67_w143, 
            w144=> c0_n67_w144, 
            w145=> c0_n67_w145, 
            w146=> c0_n67_w146, 
            w147=> c0_n67_w147, 
            w148=> c0_n67_w148, 
            w149=> c0_n67_w149, 
            w150=> c0_n67_w150, 
            w151=> c0_n67_w151, 
            w152=> c0_n67_w152, 
            w153=> c0_n67_w153, 
            w154=> c0_n67_w154, 
            w155=> c0_n67_w155, 
            w156=> c0_n67_w156, 
            w157=> c0_n67_w157, 
            w158=> c0_n67_w158, 
            w159=> c0_n67_w159, 
            w160=> c0_n67_w160, 
            w161=> c0_n67_w161, 
            w162=> c0_n67_w162, 
            w163=> c0_n67_w163, 
            w164=> c0_n67_w164, 
            w165=> c0_n67_w165, 
            w166=> c0_n67_w166, 
            w167=> c0_n67_w167, 
            w168=> c0_n67_w168, 
            w169=> c0_n67_w169, 
            w170=> c0_n67_w170, 
            w171=> c0_n67_w171, 
            w172=> c0_n67_w172, 
            w173=> c0_n67_w173, 
            w174=> c0_n67_w174, 
            w175=> c0_n67_w175, 
            w176=> c0_n67_w176, 
            w177=> c0_n67_w177, 
            w178=> c0_n67_w178, 
            w179=> c0_n67_w179, 
            w180=> c0_n67_w180, 
            w181=> c0_n67_w181, 
            w182=> c0_n67_w182, 
            w183=> c0_n67_w183, 
            w184=> c0_n67_w184, 
            w185=> c0_n67_w185, 
            w186=> c0_n67_w186, 
            w187=> c0_n67_w187, 
            w188=> c0_n67_w188, 
            w189=> c0_n67_w189, 
            w190=> c0_n67_w190, 
            w191=> c0_n67_w191, 
            w192=> c0_n67_w192, 
            w193=> c0_n67_w193, 
            w194=> c0_n67_w194, 
            w195=> c0_n67_w195, 
            w196=> c0_n67_w196, 
            w197=> c0_n67_w197, 
            w198=> c0_n67_w198, 
            w199=> c0_n67_w199, 
            w200=> c0_n67_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n67_y
   );           
            
neuron_inst_68: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n68_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n68_w1, 
            w2=> c0_n68_w2, 
            w3=> c0_n68_w3, 
            w4=> c0_n68_w4, 
            w5=> c0_n68_w5, 
            w6=> c0_n68_w6, 
            w7=> c0_n68_w7, 
            w8=> c0_n68_w8, 
            w9=> c0_n68_w9, 
            w10=> c0_n68_w10, 
            w11=> c0_n68_w11, 
            w12=> c0_n68_w12, 
            w13=> c0_n68_w13, 
            w14=> c0_n68_w14, 
            w15=> c0_n68_w15, 
            w16=> c0_n68_w16, 
            w17=> c0_n68_w17, 
            w18=> c0_n68_w18, 
            w19=> c0_n68_w19, 
            w20=> c0_n68_w20, 
            w21=> c0_n68_w21, 
            w22=> c0_n68_w22, 
            w23=> c0_n68_w23, 
            w24=> c0_n68_w24, 
            w25=> c0_n68_w25, 
            w26=> c0_n68_w26, 
            w27=> c0_n68_w27, 
            w28=> c0_n68_w28, 
            w29=> c0_n68_w29, 
            w30=> c0_n68_w30, 
            w31=> c0_n68_w31, 
            w32=> c0_n68_w32, 
            w33=> c0_n68_w33, 
            w34=> c0_n68_w34, 
            w35=> c0_n68_w35, 
            w36=> c0_n68_w36, 
            w37=> c0_n68_w37, 
            w38=> c0_n68_w38, 
            w39=> c0_n68_w39, 
            w40=> c0_n68_w40, 
            w41=> c0_n68_w41, 
            w42=> c0_n68_w42, 
            w43=> c0_n68_w43, 
            w44=> c0_n68_w44, 
            w45=> c0_n68_w45, 
            w46=> c0_n68_w46, 
            w47=> c0_n68_w47, 
            w48=> c0_n68_w48, 
            w49=> c0_n68_w49, 
            w50=> c0_n68_w50, 
            w51=> c0_n68_w51, 
            w52=> c0_n68_w52, 
            w53=> c0_n68_w53, 
            w54=> c0_n68_w54, 
            w55=> c0_n68_w55, 
            w56=> c0_n68_w56, 
            w57=> c0_n68_w57, 
            w58=> c0_n68_w58, 
            w59=> c0_n68_w59, 
            w60=> c0_n68_w60, 
            w61=> c0_n68_w61, 
            w62=> c0_n68_w62, 
            w63=> c0_n68_w63, 
            w64=> c0_n68_w64, 
            w65=> c0_n68_w65, 
            w66=> c0_n68_w66, 
            w67=> c0_n68_w67, 
            w68=> c0_n68_w68, 
            w69=> c0_n68_w69, 
            w70=> c0_n68_w70, 
            w71=> c0_n68_w71, 
            w72=> c0_n68_w72, 
            w73=> c0_n68_w73, 
            w74=> c0_n68_w74, 
            w75=> c0_n68_w75, 
            w76=> c0_n68_w76, 
            w77=> c0_n68_w77, 
            w78=> c0_n68_w78, 
            w79=> c0_n68_w79, 
            w80=> c0_n68_w80, 
            w81=> c0_n68_w81, 
            w82=> c0_n68_w82, 
            w83=> c0_n68_w83, 
            w84=> c0_n68_w84, 
            w85=> c0_n68_w85, 
            w86=> c0_n68_w86, 
            w87=> c0_n68_w87, 
            w88=> c0_n68_w88, 
            w89=> c0_n68_w89, 
            w90=> c0_n68_w90, 
            w91=> c0_n68_w91, 
            w92=> c0_n68_w92, 
            w93=> c0_n68_w93, 
            w94=> c0_n68_w94, 
            w95=> c0_n68_w95, 
            w96=> c0_n68_w96, 
            w97=> c0_n68_w97, 
            w98=> c0_n68_w98, 
            w99=> c0_n68_w99, 
            w100=> c0_n68_w100, 
            w101=> c0_n68_w101, 
            w102=> c0_n68_w102, 
            w103=> c0_n68_w103, 
            w104=> c0_n68_w104, 
            w105=> c0_n68_w105, 
            w106=> c0_n68_w106, 
            w107=> c0_n68_w107, 
            w108=> c0_n68_w108, 
            w109=> c0_n68_w109, 
            w110=> c0_n68_w110, 
            w111=> c0_n68_w111, 
            w112=> c0_n68_w112, 
            w113=> c0_n68_w113, 
            w114=> c0_n68_w114, 
            w115=> c0_n68_w115, 
            w116=> c0_n68_w116, 
            w117=> c0_n68_w117, 
            w118=> c0_n68_w118, 
            w119=> c0_n68_w119, 
            w120=> c0_n68_w120, 
            w121=> c0_n68_w121, 
            w122=> c0_n68_w122, 
            w123=> c0_n68_w123, 
            w124=> c0_n68_w124, 
            w125=> c0_n68_w125, 
            w126=> c0_n68_w126, 
            w127=> c0_n68_w127, 
            w128=> c0_n68_w128, 
            w129=> c0_n68_w129, 
            w130=> c0_n68_w130, 
            w131=> c0_n68_w131, 
            w132=> c0_n68_w132, 
            w133=> c0_n68_w133, 
            w134=> c0_n68_w134, 
            w135=> c0_n68_w135, 
            w136=> c0_n68_w136, 
            w137=> c0_n68_w137, 
            w138=> c0_n68_w138, 
            w139=> c0_n68_w139, 
            w140=> c0_n68_w140, 
            w141=> c0_n68_w141, 
            w142=> c0_n68_w142, 
            w143=> c0_n68_w143, 
            w144=> c0_n68_w144, 
            w145=> c0_n68_w145, 
            w146=> c0_n68_w146, 
            w147=> c0_n68_w147, 
            w148=> c0_n68_w148, 
            w149=> c0_n68_w149, 
            w150=> c0_n68_w150, 
            w151=> c0_n68_w151, 
            w152=> c0_n68_w152, 
            w153=> c0_n68_w153, 
            w154=> c0_n68_w154, 
            w155=> c0_n68_w155, 
            w156=> c0_n68_w156, 
            w157=> c0_n68_w157, 
            w158=> c0_n68_w158, 
            w159=> c0_n68_w159, 
            w160=> c0_n68_w160, 
            w161=> c0_n68_w161, 
            w162=> c0_n68_w162, 
            w163=> c0_n68_w163, 
            w164=> c0_n68_w164, 
            w165=> c0_n68_w165, 
            w166=> c0_n68_w166, 
            w167=> c0_n68_w167, 
            w168=> c0_n68_w168, 
            w169=> c0_n68_w169, 
            w170=> c0_n68_w170, 
            w171=> c0_n68_w171, 
            w172=> c0_n68_w172, 
            w173=> c0_n68_w173, 
            w174=> c0_n68_w174, 
            w175=> c0_n68_w175, 
            w176=> c0_n68_w176, 
            w177=> c0_n68_w177, 
            w178=> c0_n68_w178, 
            w179=> c0_n68_w179, 
            w180=> c0_n68_w180, 
            w181=> c0_n68_w181, 
            w182=> c0_n68_w182, 
            w183=> c0_n68_w183, 
            w184=> c0_n68_w184, 
            w185=> c0_n68_w185, 
            w186=> c0_n68_w186, 
            w187=> c0_n68_w187, 
            w188=> c0_n68_w188, 
            w189=> c0_n68_w189, 
            w190=> c0_n68_w190, 
            w191=> c0_n68_w191, 
            w192=> c0_n68_w192, 
            w193=> c0_n68_w193, 
            w194=> c0_n68_w194, 
            w195=> c0_n68_w195, 
            w196=> c0_n68_w196, 
            w197=> c0_n68_w197, 
            w198=> c0_n68_w198, 
            w199=> c0_n68_w199, 
            w200=> c0_n68_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n68_y
   );           
            
neuron_inst_69: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n69_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n69_w1, 
            w2=> c0_n69_w2, 
            w3=> c0_n69_w3, 
            w4=> c0_n69_w4, 
            w5=> c0_n69_w5, 
            w6=> c0_n69_w6, 
            w7=> c0_n69_w7, 
            w8=> c0_n69_w8, 
            w9=> c0_n69_w9, 
            w10=> c0_n69_w10, 
            w11=> c0_n69_w11, 
            w12=> c0_n69_w12, 
            w13=> c0_n69_w13, 
            w14=> c0_n69_w14, 
            w15=> c0_n69_w15, 
            w16=> c0_n69_w16, 
            w17=> c0_n69_w17, 
            w18=> c0_n69_w18, 
            w19=> c0_n69_w19, 
            w20=> c0_n69_w20, 
            w21=> c0_n69_w21, 
            w22=> c0_n69_w22, 
            w23=> c0_n69_w23, 
            w24=> c0_n69_w24, 
            w25=> c0_n69_w25, 
            w26=> c0_n69_w26, 
            w27=> c0_n69_w27, 
            w28=> c0_n69_w28, 
            w29=> c0_n69_w29, 
            w30=> c0_n69_w30, 
            w31=> c0_n69_w31, 
            w32=> c0_n69_w32, 
            w33=> c0_n69_w33, 
            w34=> c0_n69_w34, 
            w35=> c0_n69_w35, 
            w36=> c0_n69_w36, 
            w37=> c0_n69_w37, 
            w38=> c0_n69_w38, 
            w39=> c0_n69_w39, 
            w40=> c0_n69_w40, 
            w41=> c0_n69_w41, 
            w42=> c0_n69_w42, 
            w43=> c0_n69_w43, 
            w44=> c0_n69_w44, 
            w45=> c0_n69_w45, 
            w46=> c0_n69_w46, 
            w47=> c0_n69_w47, 
            w48=> c0_n69_w48, 
            w49=> c0_n69_w49, 
            w50=> c0_n69_w50, 
            w51=> c0_n69_w51, 
            w52=> c0_n69_w52, 
            w53=> c0_n69_w53, 
            w54=> c0_n69_w54, 
            w55=> c0_n69_w55, 
            w56=> c0_n69_w56, 
            w57=> c0_n69_w57, 
            w58=> c0_n69_w58, 
            w59=> c0_n69_w59, 
            w60=> c0_n69_w60, 
            w61=> c0_n69_w61, 
            w62=> c0_n69_w62, 
            w63=> c0_n69_w63, 
            w64=> c0_n69_w64, 
            w65=> c0_n69_w65, 
            w66=> c0_n69_w66, 
            w67=> c0_n69_w67, 
            w68=> c0_n69_w68, 
            w69=> c0_n69_w69, 
            w70=> c0_n69_w70, 
            w71=> c0_n69_w71, 
            w72=> c0_n69_w72, 
            w73=> c0_n69_w73, 
            w74=> c0_n69_w74, 
            w75=> c0_n69_w75, 
            w76=> c0_n69_w76, 
            w77=> c0_n69_w77, 
            w78=> c0_n69_w78, 
            w79=> c0_n69_w79, 
            w80=> c0_n69_w80, 
            w81=> c0_n69_w81, 
            w82=> c0_n69_w82, 
            w83=> c0_n69_w83, 
            w84=> c0_n69_w84, 
            w85=> c0_n69_w85, 
            w86=> c0_n69_w86, 
            w87=> c0_n69_w87, 
            w88=> c0_n69_w88, 
            w89=> c0_n69_w89, 
            w90=> c0_n69_w90, 
            w91=> c0_n69_w91, 
            w92=> c0_n69_w92, 
            w93=> c0_n69_w93, 
            w94=> c0_n69_w94, 
            w95=> c0_n69_w95, 
            w96=> c0_n69_w96, 
            w97=> c0_n69_w97, 
            w98=> c0_n69_w98, 
            w99=> c0_n69_w99, 
            w100=> c0_n69_w100, 
            w101=> c0_n69_w101, 
            w102=> c0_n69_w102, 
            w103=> c0_n69_w103, 
            w104=> c0_n69_w104, 
            w105=> c0_n69_w105, 
            w106=> c0_n69_w106, 
            w107=> c0_n69_w107, 
            w108=> c0_n69_w108, 
            w109=> c0_n69_w109, 
            w110=> c0_n69_w110, 
            w111=> c0_n69_w111, 
            w112=> c0_n69_w112, 
            w113=> c0_n69_w113, 
            w114=> c0_n69_w114, 
            w115=> c0_n69_w115, 
            w116=> c0_n69_w116, 
            w117=> c0_n69_w117, 
            w118=> c0_n69_w118, 
            w119=> c0_n69_w119, 
            w120=> c0_n69_w120, 
            w121=> c0_n69_w121, 
            w122=> c0_n69_w122, 
            w123=> c0_n69_w123, 
            w124=> c0_n69_w124, 
            w125=> c0_n69_w125, 
            w126=> c0_n69_w126, 
            w127=> c0_n69_w127, 
            w128=> c0_n69_w128, 
            w129=> c0_n69_w129, 
            w130=> c0_n69_w130, 
            w131=> c0_n69_w131, 
            w132=> c0_n69_w132, 
            w133=> c0_n69_w133, 
            w134=> c0_n69_w134, 
            w135=> c0_n69_w135, 
            w136=> c0_n69_w136, 
            w137=> c0_n69_w137, 
            w138=> c0_n69_w138, 
            w139=> c0_n69_w139, 
            w140=> c0_n69_w140, 
            w141=> c0_n69_w141, 
            w142=> c0_n69_w142, 
            w143=> c0_n69_w143, 
            w144=> c0_n69_w144, 
            w145=> c0_n69_w145, 
            w146=> c0_n69_w146, 
            w147=> c0_n69_w147, 
            w148=> c0_n69_w148, 
            w149=> c0_n69_w149, 
            w150=> c0_n69_w150, 
            w151=> c0_n69_w151, 
            w152=> c0_n69_w152, 
            w153=> c0_n69_w153, 
            w154=> c0_n69_w154, 
            w155=> c0_n69_w155, 
            w156=> c0_n69_w156, 
            w157=> c0_n69_w157, 
            w158=> c0_n69_w158, 
            w159=> c0_n69_w159, 
            w160=> c0_n69_w160, 
            w161=> c0_n69_w161, 
            w162=> c0_n69_w162, 
            w163=> c0_n69_w163, 
            w164=> c0_n69_w164, 
            w165=> c0_n69_w165, 
            w166=> c0_n69_w166, 
            w167=> c0_n69_w167, 
            w168=> c0_n69_w168, 
            w169=> c0_n69_w169, 
            w170=> c0_n69_w170, 
            w171=> c0_n69_w171, 
            w172=> c0_n69_w172, 
            w173=> c0_n69_w173, 
            w174=> c0_n69_w174, 
            w175=> c0_n69_w175, 
            w176=> c0_n69_w176, 
            w177=> c0_n69_w177, 
            w178=> c0_n69_w178, 
            w179=> c0_n69_w179, 
            w180=> c0_n69_w180, 
            w181=> c0_n69_w181, 
            w182=> c0_n69_w182, 
            w183=> c0_n69_w183, 
            w184=> c0_n69_w184, 
            w185=> c0_n69_w185, 
            w186=> c0_n69_w186, 
            w187=> c0_n69_w187, 
            w188=> c0_n69_w188, 
            w189=> c0_n69_w189, 
            w190=> c0_n69_w190, 
            w191=> c0_n69_w191, 
            w192=> c0_n69_w192, 
            w193=> c0_n69_w193, 
            w194=> c0_n69_w194, 
            w195=> c0_n69_w195, 
            w196=> c0_n69_w196, 
            w197=> c0_n69_w197, 
            w198=> c0_n69_w198, 
            w199=> c0_n69_w199, 
            w200=> c0_n69_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n69_y
   );           
            
neuron_inst_70: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n70_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n70_w1, 
            w2=> c0_n70_w2, 
            w3=> c0_n70_w3, 
            w4=> c0_n70_w4, 
            w5=> c0_n70_w5, 
            w6=> c0_n70_w6, 
            w7=> c0_n70_w7, 
            w8=> c0_n70_w8, 
            w9=> c0_n70_w9, 
            w10=> c0_n70_w10, 
            w11=> c0_n70_w11, 
            w12=> c0_n70_w12, 
            w13=> c0_n70_w13, 
            w14=> c0_n70_w14, 
            w15=> c0_n70_w15, 
            w16=> c0_n70_w16, 
            w17=> c0_n70_w17, 
            w18=> c0_n70_w18, 
            w19=> c0_n70_w19, 
            w20=> c0_n70_w20, 
            w21=> c0_n70_w21, 
            w22=> c0_n70_w22, 
            w23=> c0_n70_w23, 
            w24=> c0_n70_w24, 
            w25=> c0_n70_w25, 
            w26=> c0_n70_w26, 
            w27=> c0_n70_w27, 
            w28=> c0_n70_w28, 
            w29=> c0_n70_w29, 
            w30=> c0_n70_w30, 
            w31=> c0_n70_w31, 
            w32=> c0_n70_w32, 
            w33=> c0_n70_w33, 
            w34=> c0_n70_w34, 
            w35=> c0_n70_w35, 
            w36=> c0_n70_w36, 
            w37=> c0_n70_w37, 
            w38=> c0_n70_w38, 
            w39=> c0_n70_w39, 
            w40=> c0_n70_w40, 
            w41=> c0_n70_w41, 
            w42=> c0_n70_w42, 
            w43=> c0_n70_w43, 
            w44=> c0_n70_w44, 
            w45=> c0_n70_w45, 
            w46=> c0_n70_w46, 
            w47=> c0_n70_w47, 
            w48=> c0_n70_w48, 
            w49=> c0_n70_w49, 
            w50=> c0_n70_w50, 
            w51=> c0_n70_w51, 
            w52=> c0_n70_w52, 
            w53=> c0_n70_w53, 
            w54=> c0_n70_w54, 
            w55=> c0_n70_w55, 
            w56=> c0_n70_w56, 
            w57=> c0_n70_w57, 
            w58=> c0_n70_w58, 
            w59=> c0_n70_w59, 
            w60=> c0_n70_w60, 
            w61=> c0_n70_w61, 
            w62=> c0_n70_w62, 
            w63=> c0_n70_w63, 
            w64=> c0_n70_w64, 
            w65=> c0_n70_w65, 
            w66=> c0_n70_w66, 
            w67=> c0_n70_w67, 
            w68=> c0_n70_w68, 
            w69=> c0_n70_w69, 
            w70=> c0_n70_w70, 
            w71=> c0_n70_w71, 
            w72=> c0_n70_w72, 
            w73=> c0_n70_w73, 
            w74=> c0_n70_w74, 
            w75=> c0_n70_w75, 
            w76=> c0_n70_w76, 
            w77=> c0_n70_w77, 
            w78=> c0_n70_w78, 
            w79=> c0_n70_w79, 
            w80=> c0_n70_w80, 
            w81=> c0_n70_w81, 
            w82=> c0_n70_w82, 
            w83=> c0_n70_w83, 
            w84=> c0_n70_w84, 
            w85=> c0_n70_w85, 
            w86=> c0_n70_w86, 
            w87=> c0_n70_w87, 
            w88=> c0_n70_w88, 
            w89=> c0_n70_w89, 
            w90=> c0_n70_w90, 
            w91=> c0_n70_w91, 
            w92=> c0_n70_w92, 
            w93=> c0_n70_w93, 
            w94=> c0_n70_w94, 
            w95=> c0_n70_w95, 
            w96=> c0_n70_w96, 
            w97=> c0_n70_w97, 
            w98=> c0_n70_w98, 
            w99=> c0_n70_w99, 
            w100=> c0_n70_w100, 
            w101=> c0_n70_w101, 
            w102=> c0_n70_w102, 
            w103=> c0_n70_w103, 
            w104=> c0_n70_w104, 
            w105=> c0_n70_w105, 
            w106=> c0_n70_w106, 
            w107=> c0_n70_w107, 
            w108=> c0_n70_w108, 
            w109=> c0_n70_w109, 
            w110=> c0_n70_w110, 
            w111=> c0_n70_w111, 
            w112=> c0_n70_w112, 
            w113=> c0_n70_w113, 
            w114=> c0_n70_w114, 
            w115=> c0_n70_w115, 
            w116=> c0_n70_w116, 
            w117=> c0_n70_w117, 
            w118=> c0_n70_w118, 
            w119=> c0_n70_w119, 
            w120=> c0_n70_w120, 
            w121=> c0_n70_w121, 
            w122=> c0_n70_w122, 
            w123=> c0_n70_w123, 
            w124=> c0_n70_w124, 
            w125=> c0_n70_w125, 
            w126=> c0_n70_w126, 
            w127=> c0_n70_w127, 
            w128=> c0_n70_w128, 
            w129=> c0_n70_w129, 
            w130=> c0_n70_w130, 
            w131=> c0_n70_w131, 
            w132=> c0_n70_w132, 
            w133=> c0_n70_w133, 
            w134=> c0_n70_w134, 
            w135=> c0_n70_w135, 
            w136=> c0_n70_w136, 
            w137=> c0_n70_w137, 
            w138=> c0_n70_w138, 
            w139=> c0_n70_w139, 
            w140=> c0_n70_w140, 
            w141=> c0_n70_w141, 
            w142=> c0_n70_w142, 
            w143=> c0_n70_w143, 
            w144=> c0_n70_w144, 
            w145=> c0_n70_w145, 
            w146=> c0_n70_w146, 
            w147=> c0_n70_w147, 
            w148=> c0_n70_w148, 
            w149=> c0_n70_w149, 
            w150=> c0_n70_w150, 
            w151=> c0_n70_w151, 
            w152=> c0_n70_w152, 
            w153=> c0_n70_w153, 
            w154=> c0_n70_w154, 
            w155=> c0_n70_w155, 
            w156=> c0_n70_w156, 
            w157=> c0_n70_w157, 
            w158=> c0_n70_w158, 
            w159=> c0_n70_w159, 
            w160=> c0_n70_w160, 
            w161=> c0_n70_w161, 
            w162=> c0_n70_w162, 
            w163=> c0_n70_w163, 
            w164=> c0_n70_w164, 
            w165=> c0_n70_w165, 
            w166=> c0_n70_w166, 
            w167=> c0_n70_w167, 
            w168=> c0_n70_w168, 
            w169=> c0_n70_w169, 
            w170=> c0_n70_w170, 
            w171=> c0_n70_w171, 
            w172=> c0_n70_w172, 
            w173=> c0_n70_w173, 
            w174=> c0_n70_w174, 
            w175=> c0_n70_w175, 
            w176=> c0_n70_w176, 
            w177=> c0_n70_w177, 
            w178=> c0_n70_w178, 
            w179=> c0_n70_w179, 
            w180=> c0_n70_w180, 
            w181=> c0_n70_w181, 
            w182=> c0_n70_w182, 
            w183=> c0_n70_w183, 
            w184=> c0_n70_w184, 
            w185=> c0_n70_w185, 
            w186=> c0_n70_w186, 
            w187=> c0_n70_w187, 
            w188=> c0_n70_w188, 
            w189=> c0_n70_w189, 
            w190=> c0_n70_w190, 
            w191=> c0_n70_w191, 
            w192=> c0_n70_w192, 
            w193=> c0_n70_w193, 
            w194=> c0_n70_w194, 
            w195=> c0_n70_w195, 
            w196=> c0_n70_w196, 
            w197=> c0_n70_w197, 
            w198=> c0_n70_w198, 
            w199=> c0_n70_w199, 
            w200=> c0_n70_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n70_y
   );           
            
neuron_inst_71: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n71_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n71_w1, 
            w2=> c0_n71_w2, 
            w3=> c0_n71_w3, 
            w4=> c0_n71_w4, 
            w5=> c0_n71_w5, 
            w6=> c0_n71_w6, 
            w7=> c0_n71_w7, 
            w8=> c0_n71_w8, 
            w9=> c0_n71_w9, 
            w10=> c0_n71_w10, 
            w11=> c0_n71_w11, 
            w12=> c0_n71_w12, 
            w13=> c0_n71_w13, 
            w14=> c0_n71_w14, 
            w15=> c0_n71_w15, 
            w16=> c0_n71_w16, 
            w17=> c0_n71_w17, 
            w18=> c0_n71_w18, 
            w19=> c0_n71_w19, 
            w20=> c0_n71_w20, 
            w21=> c0_n71_w21, 
            w22=> c0_n71_w22, 
            w23=> c0_n71_w23, 
            w24=> c0_n71_w24, 
            w25=> c0_n71_w25, 
            w26=> c0_n71_w26, 
            w27=> c0_n71_w27, 
            w28=> c0_n71_w28, 
            w29=> c0_n71_w29, 
            w30=> c0_n71_w30, 
            w31=> c0_n71_w31, 
            w32=> c0_n71_w32, 
            w33=> c0_n71_w33, 
            w34=> c0_n71_w34, 
            w35=> c0_n71_w35, 
            w36=> c0_n71_w36, 
            w37=> c0_n71_w37, 
            w38=> c0_n71_w38, 
            w39=> c0_n71_w39, 
            w40=> c0_n71_w40, 
            w41=> c0_n71_w41, 
            w42=> c0_n71_w42, 
            w43=> c0_n71_w43, 
            w44=> c0_n71_w44, 
            w45=> c0_n71_w45, 
            w46=> c0_n71_w46, 
            w47=> c0_n71_w47, 
            w48=> c0_n71_w48, 
            w49=> c0_n71_w49, 
            w50=> c0_n71_w50, 
            w51=> c0_n71_w51, 
            w52=> c0_n71_w52, 
            w53=> c0_n71_w53, 
            w54=> c0_n71_w54, 
            w55=> c0_n71_w55, 
            w56=> c0_n71_w56, 
            w57=> c0_n71_w57, 
            w58=> c0_n71_w58, 
            w59=> c0_n71_w59, 
            w60=> c0_n71_w60, 
            w61=> c0_n71_w61, 
            w62=> c0_n71_w62, 
            w63=> c0_n71_w63, 
            w64=> c0_n71_w64, 
            w65=> c0_n71_w65, 
            w66=> c0_n71_w66, 
            w67=> c0_n71_w67, 
            w68=> c0_n71_w68, 
            w69=> c0_n71_w69, 
            w70=> c0_n71_w70, 
            w71=> c0_n71_w71, 
            w72=> c0_n71_w72, 
            w73=> c0_n71_w73, 
            w74=> c0_n71_w74, 
            w75=> c0_n71_w75, 
            w76=> c0_n71_w76, 
            w77=> c0_n71_w77, 
            w78=> c0_n71_w78, 
            w79=> c0_n71_w79, 
            w80=> c0_n71_w80, 
            w81=> c0_n71_w81, 
            w82=> c0_n71_w82, 
            w83=> c0_n71_w83, 
            w84=> c0_n71_w84, 
            w85=> c0_n71_w85, 
            w86=> c0_n71_w86, 
            w87=> c0_n71_w87, 
            w88=> c0_n71_w88, 
            w89=> c0_n71_w89, 
            w90=> c0_n71_w90, 
            w91=> c0_n71_w91, 
            w92=> c0_n71_w92, 
            w93=> c0_n71_w93, 
            w94=> c0_n71_w94, 
            w95=> c0_n71_w95, 
            w96=> c0_n71_w96, 
            w97=> c0_n71_w97, 
            w98=> c0_n71_w98, 
            w99=> c0_n71_w99, 
            w100=> c0_n71_w100, 
            w101=> c0_n71_w101, 
            w102=> c0_n71_w102, 
            w103=> c0_n71_w103, 
            w104=> c0_n71_w104, 
            w105=> c0_n71_w105, 
            w106=> c0_n71_w106, 
            w107=> c0_n71_w107, 
            w108=> c0_n71_w108, 
            w109=> c0_n71_w109, 
            w110=> c0_n71_w110, 
            w111=> c0_n71_w111, 
            w112=> c0_n71_w112, 
            w113=> c0_n71_w113, 
            w114=> c0_n71_w114, 
            w115=> c0_n71_w115, 
            w116=> c0_n71_w116, 
            w117=> c0_n71_w117, 
            w118=> c0_n71_w118, 
            w119=> c0_n71_w119, 
            w120=> c0_n71_w120, 
            w121=> c0_n71_w121, 
            w122=> c0_n71_w122, 
            w123=> c0_n71_w123, 
            w124=> c0_n71_w124, 
            w125=> c0_n71_w125, 
            w126=> c0_n71_w126, 
            w127=> c0_n71_w127, 
            w128=> c0_n71_w128, 
            w129=> c0_n71_w129, 
            w130=> c0_n71_w130, 
            w131=> c0_n71_w131, 
            w132=> c0_n71_w132, 
            w133=> c0_n71_w133, 
            w134=> c0_n71_w134, 
            w135=> c0_n71_w135, 
            w136=> c0_n71_w136, 
            w137=> c0_n71_w137, 
            w138=> c0_n71_w138, 
            w139=> c0_n71_w139, 
            w140=> c0_n71_w140, 
            w141=> c0_n71_w141, 
            w142=> c0_n71_w142, 
            w143=> c0_n71_w143, 
            w144=> c0_n71_w144, 
            w145=> c0_n71_w145, 
            w146=> c0_n71_w146, 
            w147=> c0_n71_w147, 
            w148=> c0_n71_w148, 
            w149=> c0_n71_w149, 
            w150=> c0_n71_w150, 
            w151=> c0_n71_w151, 
            w152=> c0_n71_w152, 
            w153=> c0_n71_w153, 
            w154=> c0_n71_w154, 
            w155=> c0_n71_w155, 
            w156=> c0_n71_w156, 
            w157=> c0_n71_w157, 
            w158=> c0_n71_w158, 
            w159=> c0_n71_w159, 
            w160=> c0_n71_w160, 
            w161=> c0_n71_w161, 
            w162=> c0_n71_w162, 
            w163=> c0_n71_w163, 
            w164=> c0_n71_w164, 
            w165=> c0_n71_w165, 
            w166=> c0_n71_w166, 
            w167=> c0_n71_w167, 
            w168=> c0_n71_w168, 
            w169=> c0_n71_w169, 
            w170=> c0_n71_w170, 
            w171=> c0_n71_w171, 
            w172=> c0_n71_w172, 
            w173=> c0_n71_w173, 
            w174=> c0_n71_w174, 
            w175=> c0_n71_w175, 
            w176=> c0_n71_w176, 
            w177=> c0_n71_w177, 
            w178=> c0_n71_w178, 
            w179=> c0_n71_w179, 
            w180=> c0_n71_w180, 
            w181=> c0_n71_w181, 
            w182=> c0_n71_w182, 
            w183=> c0_n71_w183, 
            w184=> c0_n71_w184, 
            w185=> c0_n71_w185, 
            w186=> c0_n71_w186, 
            w187=> c0_n71_w187, 
            w188=> c0_n71_w188, 
            w189=> c0_n71_w189, 
            w190=> c0_n71_w190, 
            w191=> c0_n71_w191, 
            w192=> c0_n71_w192, 
            w193=> c0_n71_w193, 
            w194=> c0_n71_w194, 
            w195=> c0_n71_w195, 
            w196=> c0_n71_w196, 
            w197=> c0_n71_w197, 
            w198=> c0_n71_w198, 
            w199=> c0_n71_w199, 
            w200=> c0_n71_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n71_y
   );           
            
neuron_inst_72: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n72_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n72_w1, 
            w2=> c0_n72_w2, 
            w3=> c0_n72_w3, 
            w4=> c0_n72_w4, 
            w5=> c0_n72_w5, 
            w6=> c0_n72_w6, 
            w7=> c0_n72_w7, 
            w8=> c0_n72_w8, 
            w9=> c0_n72_w9, 
            w10=> c0_n72_w10, 
            w11=> c0_n72_w11, 
            w12=> c0_n72_w12, 
            w13=> c0_n72_w13, 
            w14=> c0_n72_w14, 
            w15=> c0_n72_w15, 
            w16=> c0_n72_w16, 
            w17=> c0_n72_w17, 
            w18=> c0_n72_w18, 
            w19=> c0_n72_w19, 
            w20=> c0_n72_w20, 
            w21=> c0_n72_w21, 
            w22=> c0_n72_w22, 
            w23=> c0_n72_w23, 
            w24=> c0_n72_w24, 
            w25=> c0_n72_w25, 
            w26=> c0_n72_w26, 
            w27=> c0_n72_w27, 
            w28=> c0_n72_w28, 
            w29=> c0_n72_w29, 
            w30=> c0_n72_w30, 
            w31=> c0_n72_w31, 
            w32=> c0_n72_w32, 
            w33=> c0_n72_w33, 
            w34=> c0_n72_w34, 
            w35=> c0_n72_w35, 
            w36=> c0_n72_w36, 
            w37=> c0_n72_w37, 
            w38=> c0_n72_w38, 
            w39=> c0_n72_w39, 
            w40=> c0_n72_w40, 
            w41=> c0_n72_w41, 
            w42=> c0_n72_w42, 
            w43=> c0_n72_w43, 
            w44=> c0_n72_w44, 
            w45=> c0_n72_w45, 
            w46=> c0_n72_w46, 
            w47=> c0_n72_w47, 
            w48=> c0_n72_w48, 
            w49=> c0_n72_w49, 
            w50=> c0_n72_w50, 
            w51=> c0_n72_w51, 
            w52=> c0_n72_w52, 
            w53=> c0_n72_w53, 
            w54=> c0_n72_w54, 
            w55=> c0_n72_w55, 
            w56=> c0_n72_w56, 
            w57=> c0_n72_w57, 
            w58=> c0_n72_w58, 
            w59=> c0_n72_w59, 
            w60=> c0_n72_w60, 
            w61=> c0_n72_w61, 
            w62=> c0_n72_w62, 
            w63=> c0_n72_w63, 
            w64=> c0_n72_w64, 
            w65=> c0_n72_w65, 
            w66=> c0_n72_w66, 
            w67=> c0_n72_w67, 
            w68=> c0_n72_w68, 
            w69=> c0_n72_w69, 
            w70=> c0_n72_w70, 
            w71=> c0_n72_w71, 
            w72=> c0_n72_w72, 
            w73=> c0_n72_w73, 
            w74=> c0_n72_w74, 
            w75=> c0_n72_w75, 
            w76=> c0_n72_w76, 
            w77=> c0_n72_w77, 
            w78=> c0_n72_w78, 
            w79=> c0_n72_w79, 
            w80=> c0_n72_w80, 
            w81=> c0_n72_w81, 
            w82=> c0_n72_w82, 
            w83=> c0_n72_w83, 
            w84=> c0_n72_w84, 
            w85=> c0_n72_w85, 
            w86=> c0_n72_w86, 
            w87=> c0_n72_w87, 
            w88=> c0_n72_w88, 
            w89=> c0_n72_w89, 
            w90=> c0_n72_w90, 
            w91=> c0_n72_w91, 
            w92=> c0_n72_w92, 
            w93=> c0_n72_w93, 
            w94=> c0_n72_w94, 
            w95=> c0_n72_w95, 
            w96=> c0_n72_w96, 
            w97=> c0_n72_w97, 
            w98=> c0_n72_w98, 
            w99=> c0_n72_w99, 
            w100=> c0_n72_w100, 
            w101=> c0_n72_w101, 
            w102=> c0_n72_w102, 
            w103=> c0_n72_w103, 
            w104=> c0_n72_w104, 
            w105=> c0_n72_w105, 
            w106=> c0_n72_w106, 
            w107=> c0_n72_w107, 
            w108=> c0_n72_w108, 
            w109=> c0_n72_w109, 
            w110=> c0_n72_w110, 
            w111=> c0_n72_w111, 
            w112=> c0_n72_w112, 
            w113=> c0_n72_w113, 
            w114=> c0_n72_w114, 
            w115=> c0_n72_w115, 
            w116=> c0_n72_w116, 
            w117=> c0_n72_w117, 
            w118=> c0_n72_w118, 
            w119=> c0_n72_w119, 
            w120=> c0_n72_w120, 
            w121=> c0_n72_w121, 
            w122=> c0_n72_w122, 
            w123=> c0_n72_w123, 
            w124=> c0_n72_w124, 
            w125=> c0_n72_w125, 
            w126=> c0_n72_w126, 
            w127=> c0_n72_w127, 
            w128=> c0_n72_w128, 
            w129=> c0_n72_w129, 
            w130=> c0_n72_w130, 
            w131=> c0_n72_w131, 
            w132=> c0_n72_w132, 
            w133=> c0_n72_w133, 
            w134=> c0_n72_w134, 
            w135=> c0_n72_w135, 
            w136=> c0_n72_w136, 
            w137=> c0_n72_w137, 
            w138=> c0_n72_w138, 
            w139=> c0_n72_w139, 
            w140=> c0_n72_w140, 
            w141=> c0_n72_w141, 
            w142=> c0_n72_w142, 
            w143=> c0_n72_w143, 
            w144=> c0_n72_w144, 
            w145=> c0_n72_w145, 
            w146=> c0_n72_w146, 
            w147=> c0_n72_w147, 
            w148=> c0_n72_w148, 
            w149=> c0_n72_w149, 
            w150=> c0_n72_w150, 
            w151=> c0_n72_w151, 
            w152=> c0_n72_w152, 
            w153=> c0_n72_w153, 
            w154=> c0_n72_w154, 
            w155=> c0_n72_w155, 
            w156=> c0_n72_w156, 
            w157=> c0_n72_w157, 
            w158=> c0_n72_w158, 
            w159=> c0_n72_w159, 
            w160=> c0_n72_w160, 
            w161=> c0_n72_w161, 
            w162=> c0_n72_w162, 
            w163=> c0_n72_w163, 
            w164=> c0_n72_w164, 
            w165=> c0_n72_w165, 
            w166=> c0_n72_w166, 
            w167=> c0_n72_w167, 
            w168=> c0_n72_w168, 
            w169=> c0_n72_w169, 
            w170=> c0_n72_w170, 
            w171=> c0_n72_w171, 
            w172=> c0_n72_w172, 
            w173=> c0_n72_w173, 
            w174=> c0_n72_w174, 
            w175=> c0_n72_w175, 
            w176=> c0_n72_w176, 
            w177=> c0_n72_w177, 
            w178=> c0_n72_w178, 
            w179=> c0_n72_w179, 
            w180=> c0_n72_w180, 
            w181=> c0_n72_w181, 
            w182=> c0_n72_w182, 
            w183=> c0_n72_w183, 
            w184=> c0_n72_w184, 
            w185=> c0_n72_w185, 
            w186=> c0_n72_w186, 
            w187=> c0_n72_w187, 
            w188=> c0_n72_w188, 
            w189=> c0_n72_w189, 
            w190=> c0_n72_w190, 
            w191=> c0_n72_w191, 
            w192=> c0_n72_w192, 
            w193=> c0_n72_w193, 
            w194=> c0_n72_w194, 
            w195=> c0_n72_w195, 
            w196=> c0_n72_w196, 
            w197=> c0_n72_w197, 
            w198=> c0_n72_w198, 
            w199=> c0_n72_w199, 
            w200=> c0_n72_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n72_y
   );           
            
neuron_inst_73: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n73_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n73_w1, 
            w2=> c0_n73_w2, 
            w3=> c0_n73_w3, 
            w4=> c0_n73_w4, 
            w5=> c0_n73_w5, 
            w6=> c0_n73_w6, 
            w7=> c0_n73_w7, 
            w8=> c0_n73_w8, 
            w9=> c0_n73_w9, 
            w10=> c0_n73_w10, 
            w11=> c0_n73_w11, 
            w12=> c0_n73_w12, 
            w13=> c0_n73_w13, 
            w14=> c0_n73_w14, 
            w15=> c0_n73_w15, 
            w16=> c0_n73_w16, 
            w17=> c0_n73_w17, 
            w18=> c0_n73_w18, 
            w19=> c0_n73_w19, 
            w20=> c0_n73_w20, 
            w21=> c0_n73_w21, 
            w22=> c0_n73_w22, 
            w23=> c0_n73_w23, 
            w24=> c0_n73_w24, 
            w25=> c0_n73_w25, 
            w26=> c0_n73_w26, 
            w27=> c0_n73_w27, 
            w28=> c0_n73_w28, 
            w29=> c0_n73_w29, 
            w30=> c0_n73_w30, 
            w31=> c0_n73_w31, 
            w32=> c0_n73_w32, 
            w33=> c0_n73_w33, 
            w34=> c0_n73_w34, 
            w35=> c0_n73_w35, 
            w36=> c0_n73_w36, 
            w37=> c0_n73_w37, 
            w38=> c0_n73_w38, 
            w39=> c0_n73_w39, 
            w40=> c0_n73_w40, 
            w41=> c0_n73_w41, 
            w42=> c0_n73_w42, 
            w43=> c0_n73_w43, 
            w44=> c0_n73_w44, 
            w45=> c0_n73_w45, 
            w46=> c0_n73_w46, 
            w47=> c0_n73_w47, 
            w48=> c0_n73_w48, 
            w49=> c0_n73_w49, 
            w50=> c0_n73_w50, 
            w51=> c0_n73_w51, 
            w52=> c0_n73_w52, 
            w53=> c0_n73_w53, 
            w54=> c0_n73_w54, 
            w55=> c0_n73_w55, 
            w56=> c0_n73_w56, 
            w57=> c0_n73_w57, 
            w58=> c0_n73_w58, 
            w59=> c0_n73_w59, 
            w60=> c0_n73_w60, 
            w61=> c0_n73_w61, 
            w62=> c0_n73_w62, 
            w63=> c0_n73_w63, 
            w64=> c0_n73_w64, 
            w65=> c0_n73_w65, 
            w66=> c0_n73_w66, 
            w67=> c0_n73_w67, 
            w68=> c0_n73_w68, 
            w69=> c0_n73_w69, 
            w70=> c0_n73_w70, 
            w71=> c0_n73_w71, 
            w72=> c0_n73_w72, 
            w73=> c0_n73_w73, 
            w74=> c0_n73_w74, 
            w75=> c0_n73_w75, 
            w76=> c0_n73_w76, 
            w77=> c0_n73_w77, 
            w78=> c0_n73_w78, 
            w79=> c0_n73_w79, 
            w80=> c0_n73_w80, 
            w81=> c0_n73_w81, 
            w82=> c0_n73_w82, 
            w83=> c0_n73_w83, 
            w84=> c0_n73_w84, 
            w85=> c0_n73_w85, 
            w86=> c0_n73_w86, 
            w87=> c0_n73_w87, 
            w88=> c0_n73_w88, 
            w89=> c0_n73_w89, 
            w90=> c0_n73_w90, 
            w91=> c0_n73_w91, 
            w92=> c0_n73_w92, 
            w93=> c0_n73_w93, 
            w94=> c0_n73_w94, 
            w95=> c0_n73_w95, 
            w96=> c0_n73_w96, 
            w97=> c0_n73_w97, 
            w98=> c0_n73_w98, 
            w99=> c0_n73_w99, 
            w100=> c0_n73_w100, 
            w101=> c0_n73_w101, 
            w102=> c0_n73_w102, 
            w103=> c0_n73_w103, 
            w104=> c0_n73_w104, 
            w105=> c0_n73_w105, 
            w106=> c0_n73_w106, 
            w107=> c0_n73_w107, 
            w108=> c0_n73_w108, 
            w109=> c0_n73_w109, 
            w110=> c0_n73_w110, 
            w111=> c0_n73_w111, 
            w112=> c0_n73_w112, 
            w113=> c0_n73_w113, 
            w114=> c0_n73_w114, 
            w115=> c0_n73_w115, 
            w116=> c0_n73_w116, 
            w117=> c0_n73_w117, 
            w118=> c0_n73_w118, 
            w119=> c0_n73_w119, 
            w120=> c0_n73_w120, 
            w121=> c0_n73_w121, 
            w122=> c0_n73_w122, 
            w123=> c0_n73_w123, 
            w124=> c0_n73_w124, 
            w125=> c0_n73_w125, 
            w126=> c0_n73_w126, 
            w127=> c0_n73_w127, 
            w128=> c0_n73_w128, 
            w129=> c0_n73_w129, 
            w130=> c0_n73_w130, 
            w131=> c0_n73_w131, 
            w132=> c0_n73_w132, 
            w133=> c0_n73_w133, 
            w134=> c0_n73_w134, 
            w135=> c0_n73_w135, 
            w136=> c0_n73_w136, 
            w137=> c0_n73_w137, 
            w138=> c0_n73_w138, 
            w139=> c0_n73_w139, 
            w140=> c0_n73_w140, 
            w141=> c0_n73_w141, 
            w142=> c0_n73_w142, 
            w143=> c0_n73_w143, 
            w144=> c0_n73_w144, 
            w145=> c0_n73_w145, 
            w146=> c0_n73_w146, 
            w147=> c0_n73_w147, 
            w148=> c0_n73_w148, 
            w149=> c0_n73_w149, 
            w150=> c0_n73_w150, 
            w151=> c0_n73_w151, 
            w152=> c0_n73_w152, 
            w153=> c0_n73_w153, 
            w154=> c0_n73_w154, 
            w155=> c0_n73_w155, 
            w156=> c0_n73_w156, 
            w157=> c0_n73_w157, 
            w158=> c0_n73_w158, 
            w159=> c0_n73_w159, 
            w160=> c0_n73_w160, 
            w161=> c0_n73_w161, 
            w162=> c0_n73_w162, 
            w163=> c0_n73_w163, 
            w164=> c0_n73_w164, 
            w165=> c0_n73_w165, 
            w166=> c0_n73_w166, 
            w167=> c0_n73_w167, 
            w168=> c0_n73_w168, 
            w169=> c0_n73_w169, 
            w170=> c0_n73_w170, 
            w171=> c0_n73_w171, 
            w172=> c0_n73_w172, 
            w173=> c0_n73_w173, 
            w174=> c0_n73_w174, 
            w175=> c0_n73_w175, 
            w176=> c0_n73_w176, 
            w177=> c0_n73_w177, 
            w178=> c0_n73_w178, 
            w179=> c0_n73_w179, 
            w180=> c0_n73_w180, 
            w181=> c0_n73_w181, 
            w182=> c0_n73_w182, 
            w183=> c0_n73_w183, 
            w184=> c0_n73_w184, 
            w185=> c0_n73_w185, 
            w186=> c0_n73_w186, 
            w187=> c0_n73_w187, 
            w188=> c0_n73_w188, 
            w189=> c0_n73_w189, 
            w190=> c0_n73_w190, 
            w191=> c0_n73_w191, 
            w192=> c0_n73_w192, 
            w193=> c0_n73_w193, 
            w194=> c0_n73_w194, 
            w195=> c0_n73_w195, 
            w196=> c0_n73_w196, 
            w197=> c0_n73_w197, 
            w198=> c0_n73_w198, 
            w199=> c0_n73_w199, 
            w200=> c0_n73_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n73_y
   );           
            
neuron_inst_74: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n74_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n74_w1, 
            w2=> c0_n74_w2, 
            w3=> c0_n74_w3, 
            w4=> c0_n74_w4, 
            w5=> c0_n74_w5, 
            w6=> c0_n74_w6, 
            w7=> c0_n74_w7, 
            w8=> c0_n74_w8, 
            w9=> c0_n74_w9, 
            w10=> c0_n74_w10, 
            w11=> c0_n74_w11, 
            w12=> c0_n74_w12, 
            w13=> c0_n74_w13, 
            w14=> c0_n74_w14, 
            w15=> c0_n74_w15, 
            w16=> c0_n74_w16, 
            w17=> c0_n74_w17, 
            w18=> c0_n74_w18, 
            w19=> c0_n74_w19, 
            w20=> c0_n74_w20, 
            w21=> c0_n74_w21, 
            w22=> c0_n74_w22, 
            w23=> c0_n74_w23, 
            w24=> c0_n74_w24, 
            w25=> c0_n74_w25, 
            w26=> c0_n74_w26, 
            w27=> c0_n74_w27, 
            w28=> c0_n74_w28, 
            w29=> c0_n74_w29, 
            w30=> c0_n74_w30, 
            w31=> c0_n74_w31, 
            w32=> c0_n74_w32, 
            w33=> c0_n74_w33, 
            w34=> c0_n74_w34, 
            w35=> c0_n74_w35, 
            w36=> c0_n74_w36, 
            w37=> c0_n74_w37, 
            w38=> c0_n74_w38, 
            w39=> c0_n74_w39, 
            w40=> c0_n74_w40, 
            w41=> c0_n74_w41, 
            w42=> c0_n74_w42, 
            w43=> c0_n74_w43, 
            w44=> c0_n74_w44, 
            w45=> c0_n74_w45, 
            w46=> c0_n74_w46, 
            w47=> c0_n74_w47, 
            w48=> c0_n74_w48, 
            w49=> c0_n74_w49, 
            w50=> c0_n74_w50, 
            w51=> c0_n74_w51, 
            w52=> c0_n74_w52, 
            w53=> c0_n74_w53, 
            w54=> c0_n74_w54, 
            w55=> c0_n74_w55, 
            w56=> c0_n74_w56, 
            w57=> c0_n74_w57, 
            w58=> c0_n74_w58, 
            w59=> c0_n74_w59, 
            w60=> c0_n74_w60, 
            w61=> c0_n74_w61, 
            w62=> c0_n74_w62, 
            w63=> c0_n74_w63, 
            w64=> c0_n74_w64, 
            w65=> c0_n74_w65, 
            w66=> c0_n74_w66, 
            w67=> c0_n74_w67, 
            w68=> c0_n74_w68, 
            w69=> c0_n74_w69, 
            w70=> c0_n74_w70, 
            w71=> c0_n74_w71, 
            w72=> c0_n74_w72, 
            w73=> c0_n74_w73, 
            w74=> c0_n74_w74, 
            w75=> c0_n74_w75, 
            w76=> c0_n74_w76, 
            w77=> c0_n74_w77, 
            w78=> c0_n74_w78, 
            w79=> c0_n74_w79, 
            w80=> c0_n74_w80, 
            w81=> c0_n74_w81, 
            w82=> c0_n74_w82, 
            w83=> c0_n74_w83, 
            w84=> c0_n74_w84, 
            w85=> c0_n74_w85, 
            w86=> c0_n74_w86, 
            w87=> c0_n74_w87, 
            w88=> c0_n74_w88, 
            w89=> c0_n74_w89, 
            w90=> c0_n74_w90, 
            w91=> c0_n74_w91, 
            w92=> c0_n74_w92, 
            w93=> c0_n74_w93, 
            w94=> c0_n74_w94, 
            w95=> c0_n74_w95, 
            w96=> c0_n74_w96, 
            w97=> c0_n74_w97, 
            w98=> c0_n74_w98, 
            w99=> c0_n74_w99, 
            w100=> c0_n74_w100, 
            w101=> c0_n74_w101, 
            w102=> c0_n74_w102, 
            w103=> c0_n74_w103, 
            w104=> c0_n74_w104, 
            w105=> c0_n74_w105, 
            w106=> c0_n74_w106, 
            w107=> c0_n74_w107, 
            w108=> c0_n74_w108, 
            w109=> c0_n74_w109, 
            w110=> c0_n74_w110, 
            w111=> c0_n74_w111, 
            w112=> c0_n74_w112, 
            w113=> c0_n74_w113, 
            w114=> c0_n74_w114, 
            w115=> c0_n74_w115, 
            w116=> c0_n74_w116, 
            w117=> c0_n74_w117, 
            w118=> c0_n74_w118, 
            w119=> c0_n74_w119, 
            w120=> c0_n74_w120, 
            w121=> c0_n74_w121, 
            w122=> c0_n74_w122, 
            w123=> c0_n74_w123, 
            w124=> c0_n74_w124, 
            w125=> c0_n74_w125, 
            w126=> c0_n74_w126, 
            w127=> c0_n74_w127, 
            w128=> c0_n74_w128, 
            w129=> c0_n74_w129, 
            w130=> c0_n74_w130, 
            w131=> c0_n74_w131, 
            w132=> c0_n74_w132, 
            w133=> c0_n74_w133, 
            w134=> c0_n74_w134, 
            w135=> c0_n74_w135, 
            w136=> c0_n74_w136, 
            w137=> c0_n74_w137, 
            w138=> c0_n74_w138, 
            w139=> c0_n74_w139, 
            w140=> c0_n74_w140, 
            w141=> c0_n74_w141, 
            w142=> c0_n74_w142, 
            w143=> c0_n74_w143, 
            w144=> c0_n74_w144, 
            w145=> c0_n74_w145, 
            w146=> c0_n74_w146, 
            w147=> c0_n74_w147, 
            w148=> c0_n74_w148, 
            w149=> c0_n74_w149, 
            w150=> c0_n74_w150, 
            w151=> c0_n74_w151, 
            w152=> c0_n74_w152, 
            w153=> c0_n74_w153, 
            w154=> c0_n74_w154, 
            w155=> c0_n74_w155, 
            w156=> c0_n74_w156, 
            w157=> c0_n74_w157, 
            w158=> c0_n74_w158, 
            w159=> c0_n74_w159, 
            w160=> c0_n74_w160, 
            w161=> c0_n74_w161, 
            w162=> c0_n74_w162, 
            w163=> c0_n74_w163, 
            w164=> c0_n74_w164, 
            w165=> c0_n74_w165, 
            w166=> c0_n74_w166, 
            w167=> c0_n74_w167, 
            w168=> c0_n74_w168, 
            w169=> c0_n74_w169, 
            w170=> c0_n74_w170, 
            w171=> c0_n74_w171, 
            w172=> c0_n74_w172, 
            w173=> c0_n74_w173, 
            w174=> c0_n74_w174, 
            w175=> c0_n74_w175, 
            w176=> c0_n74_w176, 
            w177=> c0_n74_w177, 
            w178=> c0_n74_w178, 
            w179=> c0_n74_w179, 
            w180=> c0_n74_w180, 
            w181=> c0_n74_w181, 
            w182=> c0_n74_w182, 
            w183=> c0_n74_w183, 
            w184=> c0_n74_w184, 
            w185=> c0_n74_w185, 
            w186=> c0_n74_w186, 
            w187=> c0_n74_w187, 
            w188=> c0_n74_w188, 
            w189=> c0_n74_w189, 
            w190=> c0_n74_w190, 
            w191=> c0_n74_w191, 
            w192=> c0_n74_w192, 
            w193=> c0_n74_w193, 
            w194=> c0_n74_w194, 
            w195=> c0_n74_w195, 
            w196=> c0_n74_w196, 
            w197=> c0_n74_w197, 
            w198=> c0_n74_w198, 
            w199=> c0_n74_w199, 
            w200=> c0_n74_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n74_y
   );           
            
neuron_inst_75: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n75_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n75_w1, 
            w2=> c0_n75_w2, 
            w3=> c0_n75_w3, 
            w4=> c0_n75_w4, 
            w5=> c0_n75_w5, 
            w6=> c0_n75_w6, 
            w7=> c0_n75_w7, 
            w8=> c0_n75_w8, 
            w9=> c0_n75_w9, 
            w10=> c0_n75_w10, 
            w11=> c0_n75_w11, 
            w12=> c0_n75_w12, 
            w13=> c0_n75_w13, 
            w14=> c0_n75_w14, 
            w15=> c0_n75_w15, 
            w16=> c0_n75_w16, 
            w17=> c0_n75_w17, 
            w18=> c0_n75_w18, 
            w19=> c0_n75_w19, 
            w20=> c0_n75_w20, 
            w21=> c0_n75_w21, 
            w22=> c0_n75_w22, 
            w23=> c0_n75_w23, 
            w24=> c0_n75_w24, 
            w25=> c0_n75_w25, 
            w26=> c0_n75_w26, 
            w27=> c0_n75_w27, 
            w28=> c0_n75_w28, 
            w29=> c0_n75_w29, 
            w30=> c0_n75_w30, 
            w31=> c0_n75_w31, 
            w32=> c0_n75_w32, 
            w33=> c0_n75_w33, 
            w34=> c0_n75_w34, 
            w35=> c0_n75_w35, 
            w36=> c0_n75_w36, 
            w37=> c0_n75_w37, 
            w38=> c0_n75_w38, 
            w39=> c0_n75_w39, 
            w40=> c0_n75_w40, 
            w41=> c0_n75_w41, 
            w42=> c0_n75_w42, 
            w43=> c0_n75_w43, 
            w44=> c0_n75_w44, 
            w45=> c0_n75_w45, 
            w46=> c0_n75_w46, 
            w47=> c0_n75_w47, 
            w48=> c0_n75_w48, 
            w49=> c0_n75_w49, 
            w50=> c0_n75_w50, 
            w51=> c0_n75_w51, 
            w52=> c0_n75_w52, 
            w53=> c0_n75_w53, 
            w54=> c0_n75_w54, 
            w55=> c0_n75_w55, 
            w56=> c0_n75_w56, 
            w57=> c0_n75_w57, 
            w58=> c0_n75_w58, 
            w59=> c0_n75_w59, 
            w60=> c0_n75_w60, 
            w61=> c0_n75_w61, 
            w62=> c0_n75_w62, 
            w63=> c0_n75_w63, 
            w64=> c0_n75_w64, 
            w65=> c0_n75_w65, 
            w66=> c0_n75_w66, 
            w67=> c0_n75_w67, 
            w68=> c0_n75_w68, 
            w69=> c0_n75_w69, 
            w70=> c0_n75_w70, 
            w71=> c0_n75_w71, 
            w72=> c0_n75_w72, 
            w73=> c0_n75_w73, 
            w74=> c0_n75_w74, 
            w75=> c0_n75_w75, 
            w76=> c0_n75_w76, 
            w77=> c0_n75_w77, 
            w78=> c0_n75_w78, 
            w79=> c0_n75_w79, 
            w80=> c0_n75_w80, 
            w81=> c0_n75_w81, 
            w82=> c0_n75_w82, 
            w83=> c0_n75_w83, 
            w84=> c0_n75_w84, 
            w85=> c0_n75_w85, 
            w86=> c0_n75_w86, 
            w87=> c0_n75_w87, 
            w88=> c0_n75_w88, 
            w89=> c0_n75_w89, 
            w90=> c0_n75_w90, 
            w91=> c0_n75_w91, 
            w92=> c0_n75_w92, 
            w93=> c0_n75_w93, 
            w94=> c0_n75_w94, 
            w95=> c0_n75_w95, 
            w96=> c0_n75_w96, 
            w97=> c0_n75_w97, 
            w98=> c0_n75_w98, 
            w99=> c0_n75_w99, 
            w100=> c0_n75_w100, 
            w101=> c0_n75_w101, 
            w102=> c0_n75_w102, 
            w103=> c0_n75_w103, 
            w104=> c0_n75_w104, 
            w105=> c0_n75_w105, 
            w106=> c0_n75_w106, 
            w107=> c0_n75_w107, 
            w108=> c0_n75_w108, 
            w109=> c0_n75_w109, 
            w110=> c0_n75_w110, 
            w111=> c0_n75_w111, 
            w112=> c0_n75_w112, 
            w113=> c0_n75_w113, 
            w114=> c0_n75_w114, 
            w115=> c0_n75_w115, 
            w116=> c0_n75_w116, 
            w117=> c0_n75_w117, 
            w118=> c0_n75_w118, 
            w119=> c0_n75_w119, 
            w120=> c0_n75_w120, 
            w121=> c0_n75_w121, 
            w122=> c0_n75_w122, 
            w123=> c0_n75_w123, 
            w124=> c0_n75_w124, 
            w125=> c0_n75_w125, 
            w126=> c0_n75_w126, 
            w127=> c0_n75_w127, 
            w128=> c0_n75_w128, 
            w129=> c0_n75_w129, 
            w130=> c0_n75_w130, 
            w131=> c0_n75_w131, 
            w132=> c0_n75_w132, 
            w133=> c0_n75_w133, 
            w134=> c0_n75_w134, 
            w135=> c0_n75_w135, 
            w136=> c0_n75_w136, 
            w137=> c0_n75_w137, 
            w138=> c0_n75_w138, 
            w139=> c0_n75_w139, 
            w140=> c0_n75_w140, 
            w141=> c0_n75_w141, 
            w142=> c0_n75_w142, 
            w143=> c0_n75_w143, 
            w144=> c0_n75_w144, 
            w145=> c0_n75_w145, 
            w146=> c0_n75_w146, 
            w147=> c0_n75_w147, 
            w148=> c0_n75_w148, 
            w149=> c0_n75_w149, 
            w150=> c0_n75_w150, 
            w151=> c0_n75_w151, 
            w152=> c0_n75_w152, 
            w153=> c0_n75_w153, 
            w154=> c0_n75_w154, 
            w155=> c0_n75_w155, 
            w156=> c0_n75_w156, 
            w157=> c0_n75_w157, 
            w158=> c0_n75_w158, 
            w159=> c0_n75_w159, 
            w160=> c0_n75_w160, 
            w161=> c0_n75_w161, 
            w162=> c0_n75_w162, 
            w163=> c0_n75_w163, 
            w164=> c0_n75_w164, 
            w165=> c0_n75_w165, 
            w166=> c0_n75_w166, 
            w167=> c0_n75_w167, 
            w168=> c0_n75_w168, 
            w169=> c0_n75_w169, 
            w170=> c0_n75_w170, 
            w171=> c0_n75_w171, 
            w172=> c0_n75_w172, 
            w173=> c0_n75_w173, 
            w174=> c0_n75_w174, 
            w175=> c0_n75_w175, 
            w176=> c0_n75_w176, 
            w177=> c0_n75_w177, 
            w178=> c0_n75_w178, 
            w179=> c0_n75_w179, 
            w180=> c0_n75_w180, 
            w181=> c0_n75_w181, 
            w182=> c0_n75_w182, 
            w183=> c0_n75_w183, 
            w184=> c0_n75_w184, 
            w185=> c0_n75_w185, 
            w186=> c0_n75_w186, 
            w187=> c0_n75_w187, 
            w188=> c0_n75_w188, 
            w189=> c0_n75_w189, 
            w190=> c0_n75_w190, 
            w191=> c0_n75_w191, 
            w192=> c0_n75_w192, 
            w193=> c0_n75_w193, 
            w194=> c0_n75_w194, 
            w195=> c0_n75_w195, 
            w196=> c0_n75_w196, 
            w197=> c0_n75_w197, 
            w198=> c0_n75_w198, 
            w199=> c0_n75_w199, 
            w200=> c0_n75_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n75_y
   );           
            
neuron_inst_76: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n76_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n76_w1, 
            w2=> c0_n76_w2, 
            w3=> c0_n76_w3, 
            w4=> c0_n76_w4, 
            w5=> c0_n76_w5, 
            w6=> c0_n76_w6, 
            w7=> c0_n76_w7, 
            w8=> c0_n76_w8, 
            w9=> c0_n76_w9, 
            w10=> c0_n76_w10, 
            w11=> c0_n76_w11, 
            w12=> c0_n76_w12, 
            w13=> c0_n76_w13, 
            w14=> c0_n76_w14, 
            w15=> c0_n76_w15, 
            w16=> c0_n76_w16, 
            w17=> c0_n76_w17, 
            w18=> c0_n76_w18, 
            w19=> c0_n76_w19, 
            w20=> c0_n76_w20, 
            w21=> c0_n76_w21, 
            w22=> c0_n76_w22, 
            w23=> c0_n76_w23, 
            w24=> c0_n76_w24, 
            w25=> c0_n76_w25, 
            w26=> c0_n76_w26, 
            w27=> c0_n76_w27, 
            w28=> c0_n76_w28, 
            w29=> c0_n76_w29, 
            w30=> c0_n76_w30, 
            w31=> c0_n76_w31, 
            w32=> c0_n76_w32, 
            w33=> c0_n76_w33, 
            w34=> c0_n76_w34, 
            w35=> c0_n76_w35, 
            w36=> c0_n76_w36, 
            w37=> c0_n76_w37, 
            w38=> c0_n76_w38, 
            w39=> c0_n76_w39, 
            w40=> c0_n76_w40, 
            w41=> c0_n76_w41, 
            w42=> c0_n76_w42, 
            w43=> c0_n76_w43, 
            w44=> c0_n76_w44, 
            w45=> c0_n76_w45, 
            w46=> c0_n76_w46, 
            w47=> c0_n76_w47, 
            w48=> c0_n76_w48, 
            w49=> c0_n76_w49, 
            w50=> c0_n76_w50, 
            w51=> c0_n76_w51, 
            w52=> c0_n76_w52, 
            w53=> c0_n76_w53, 
            w54=> c0_n76_w54, 
            w55=> c0_n76_w55, 
            w56=> c0_n76_w56, 
            w57=> c0_n76_w57, 
            w58=> c0_n76_w58, 
            w59=> c0_n76_w59, 
            w60=> c0_n76_w60, 
            w61=> c0_n76_w61, 
            w62=> c0_n76_w62, 
            w63=> c0_n76_w63, 
            w64=> c0_n76_w64, 
            w65=> c0_n76_w65, 
            w66=> c0_n76_w66, 
            w67=> c0_n76_w67, 
            w68=> c0_n76_w68, 
            w69=> c0_n76_w69, 
            w70=> c0_n76_w70, 
            w71=> c0_n76_w71, 
            w72=> c0_n76_w72, 
            w73=> c0_n76_w73, 
            w74=> c0_n76_w74, 
            w75=> c0_n76_w75, 
            w76=> c0_n76_w76, 
            w77=> c0_n76_w77, 
            w78=> c0_n76_w78, 
            w79=> c0_n76_w79, 
            w80=> c0_n76_w80, 
            w81=> c0_n76_w81, 
            w82=> c0_n76_w82, 
            w83=> c0_n76_w83, 
            w84=> c0_n76_w84, 
            w85=> c0_n76_w85, 
            w86=> c0_n76_w86, 
            w87=> c0_n76_w87, 
            w88=> c0_n76_w88, 
            w89=> c0_n76_w89, 
            w90=> c0_n76_w90, 
            w91=> c0_n76_w91, 
            w92=> c0_n76_w92, 
            w93=> c0_n76_w93, 
            w94=> c0_n76_w94, 
            w95=> c0_n76_w95, 
            w96=> c0_n76_w96, 
            w97=> c0_n76_w97, 
            w98=> c0_n76_w98, 
            w99=> c0_n76_w99, 
            w100=> c0_n76_w100, 
            w101=> c0_n76_w101, 
            w102=> c0_n76_w102, 
            w103=> c0_n76_w103, 
            w104=> c0_n76_w104, 
            w105=> c0_n76_w105, 
            w106=> c0_n76_w106, 
            w107=> c0_n76_w107, 
            w108=> c0_n76_w108, 
            w109=> c0_n76_w109, 
            w110=> c0_n76_w110, 
            w111=> c0_n76_w111, 
            w112=> c0_n76_w112, 
            w113=> c0_n76_w113, 
            w114=> c0_n76_w114, 
            w115=> c0_n76_w115, 
            w116=> c0_n76_w116, 
            w117=> c0_n76_w117, 
            w118=> c0_n76_w118, 
            w119=> c0_n76_w119, 
            w120=> c0_n76_w120, 
            w121=> c0_n76_w121, 
            w122=> c0_n76_w122, 
            w123=> c0_n76_w123, 
            w124=> c0_n76_w124, 
            w125=> c0_n76_w125, 
            w126=> c0_n76_w126, 
            w127=> c0_n76_w127, 
            w128=> c0_n76_w128, 
            w129=> c0_n76_w129, 
            w130=> c0_n76_w130, 
            w131=> c0_n76_w131, 
            w132=> c0_n76_w132, 
            w133=> c0_n76_w133, 
            w134=> c0_n76_w134, 
            w135=> c0_n76_w135, 
            w136=> c0_n76_w136, 
            w137=> c0_n76_w137, 
            w138=> c0_n76_w138, 
            w139=> c0_n76_w139, 
            w140=> c0_n76_w140, 
            w141=> c0_n76_w141, 
            w142=> c0_n76_w142, 
            w143=> c0_n76_w143, 
            w144=> c0_n76_w144, 
            w145=> c0_n76_w145, 
            w146=> c0_n76_w146, 
            w147=> c0_n76_w147, 
            w148=> c0_n76_w148, 
            w149=> c0_n76_w149, 
            w150=> c0_n76_w150, 
            w151=> c0_n76_w151, 
            w152=> c0_n76_w152, 
            w153=> c0_n76_w153, 
            w154=> c0_n76_w154, 
            w155=> c0_n76_w155, 
            w156=> c0_n76_w156, 
            w157=> c0_n76_w157, 
            w158=> c0_n76_w158, 
            w159=> c0_n76_w159, 
            w160=> c0_n76_w160, 
            w161=> c0_n76_w161, 
            w162=> c0_n76_w162, 
            w163=> c0_n76_w163, 
            w164=> c0_n76_w164, 
            w165=> c0_n76_w165, 
            w166=> c0_n76_w166, 
            w167=> c0_n76_w167, 
            w168=> c0_n76_w168, 
            w169=> c0_n76_w169, 
            w170=> c0_n76_w170, 
            w171=> c0_n76_w171, 
            w172=> c0_n76_w172, 
            w173=> c0_n76_w173, 
            w174=> c0_n76_w174, 
            w175=> c0_n76_w175, 
            w176=> c0_n76_w176, 
            w177=> c0_n76_w177, 
            w178=> c0_n76_w178, 
            w179=> c0_n76_w179, 
            w180=> c0_n76_w180, 
            w181=> c0_n76_w181, 
            w182=> c0_n76_w182, 
            w183=> c0_n76_w183, 
            w184=> c0_n76_w184, 
            w185=> c0_n76_w185, 
            w186=> c0_n76_w186, 
            w187=> c0_n76_w187, 
            w188=> c0_n76_w188, 
            w189=> c0_n76_w189, 
            w190=> c0_n76_w190, 
            w191=> c0_n76_w191, 
            w192=> c0_n76_w192, 
            w193=> c0_n76_w193, 
            w194=> c0_n76_w194, 
            w195=> c0_n76_w195, 
            w196=> c0_n76_w196, 
            w197=> c0_n76_w197, 
            w198=> c0_n76_w198, 
            w199=> c0_n76_w199, 
            w200=> c0_n76_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n76_y
   );           
            
neuron_inst_77: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n77_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n77_w1, 
            w2=> c0_n77_w2, 
            w3=> c0_n77_w3, 
            w4=> c0_n77_w4, 
            w5=> c0_n77_w5, 
            w6=> c0_n77_w6, 
            w7=> c0_n77_w7, 
            w8=> c0_n77_w8, 
            w9=> c0_n77_w9, 
            w10=> c0_n77_w10, 
            w11=> c0_n77_w11, 
            w12=> c0_n77_w12, 
            w13=> c0_n77_w13, 
            w14=> c0_n77_w14, 
            w15=> c0_n77_w15, 
            w16=> c0_n77_w16, 
            w17=> c0_n77_w17, 
            w18=> c0_n77_w18, 
            w19=> c0_n77_w19, 
            w20=> c0_n77_w20, 
            w21=> c0_n77_w21, 
            w22=> c0_n77_w22, 
            w23=> c0_n77_w23, 
            w24=> c0_n77_w24, 
            w25=> c0_n77_w25, 
            w26=> c0_n77_w26, 
            w27=> c0_n77_w27, 
            w28=> c0_n77_w28, 
            w29=> c0_n77_w29, 
            w30=> c0_n77_w30, 
            w31=> c0_n77_w31, 
            w32=> c0_n77_w32, 
            w33=> c0_n77_w33, 
            w34=> c0_n77_w34, 
            w35=> c0_n77_w35, 
            w36=> c0_n77_w36, 
            w37=> c0_n77_w37, 
            w38=> c0_n77_w38, 
            w39=> c0_n77_w39, 
            w40=> c0_n77_w40, 
            w41=> c0_n77_w41, 
            w42=> c0_n77_w42, 
            w43=> c0_n77_w43, 
            w44=> c0_n77_w44, 
            w45=> c0_n77_w45, 
            w46=> c0_n77_w46, 
            w47=> c0_n77_w47, 
            w48=> c0_n77_w48, 
            w49=> c0_n77_w49, 
            w50=> c0_n77_w50, 
            w51=> c0_n77_w51, 
            w52=> c0_n77_w52, 
            w53=> c0_n77_w53, 
            w54=> c0_n77_w54, 
            w55=> c0_n77_w55, 
            w56=> c0_n77_w56, 
            w57=> c0_n77_w57, 
            w58=> c0_n77_w58, 
            w59=> c0_n77_w59, 
            w60=> c0_n77_w60, 
            w61=> c0_n77_w61, 
            w62=> c0_n77_w62, 
            w63=> c0_n77_w63, 
            w64=> c0_n77_w64, 
            w65=> c0_n77_w65, 
            w66=> c0_n77_w66, 
            w67=> c0_n77_w67, 
            w68=> c0_n77_w68, 
            w69=> c0_n77_w69, 
            w70=> c0_n77_w70, 
            w71=> c0_n77_w71, 
            w72=> c0_n77_w72, 
            w73=> c0_n77_w73, 
            w74=> c0_n77_w74, 
            w75=> c0_n77_w75, 
            w76=> c0_n77_w76, 
            w77=> c0_n77_w77, 
            w78=> c0_n77_w78, 
            w79=> c0_n77_w79, 
            w80=> c0_n77_w80, 
            w81=> c0_n77_w81, 
            w82=> c0_n77_w82, 
            w83=> c0_n77_w83, 
            w84=> c0_n77_w84, 
            w85=> c0_n77_w85, 
            w86=> c0_n77_w86, 
            w87=> c0_n77_w87, 
            w88=> c0_n77_w88, 
            w89=> c0_n77_w89, 
            w90=> c0_n77_w90, 
            w91=> c0_n77_w91, 
            w92=> c0_n77_w92, 
            w93=> c0_n77_w93, 
            w94=> c0_n77_w94, 
            w95=> c0_n77_w95, 
            w96=> c0_n77_w96, 
            w97=> c0_n77_w97, 
            w98=> c0_n77_w98, 
            w99=> c0_n77_w99, 
            w100=> c0_n77_w100, 
            w101=> c0_n77_w101, 
            w102=> c0_n77_w102, 
            w103=> c0_n77_w103, 
            w104=> c0_n77_w104, 
            w105=> c0_n77_w105, 
            w106=> c0_n77_w106, 
            w107=> c0_n77_w107, 
            w108=> c0_n77_w108, 
            w109=> c0_n77_w109, 
            w110=> c0_n77_w110, 
            w111=> c0_n77_w111, 
            w112=> c0_n77_w112, 
            w113=> c0_n77_w113, 
            w114=> c0_n77_w114, 
            w115=> c0_n77_w115, 
            w116=> c0_n77_w116, 
            w117=> c0_n77_w117, 
            w118=> c0_n77_w118, 
            w119=> c0_n77_w119, 
            w120=> c0_n77_w120, 
            w121=> c0_n77_w121, 
            w122=> c0_n77_w122, 
            w123=> c0_n77_w123, 
            w124=> c0_n77_w124, 
            w125=> c0_n77_w125, 
            w126=> c0_n77_w126, 
            w127=> c0_n77_w127, 
            w128=> c0_n77_w128, 
            w129=> c0_n77_w129, 
            w130=> c0_n77_w130, 
            w131=> c0_n77_w131, 
            w132=> c0_n77_w132, 
            w133=> c0_n77_w133, 
            w134=> c0_n77_w134, 
            w135=> c0_n77_w135, 
            w136=> c0_n77_w136, 
            w137=> c0_n77_w137, 
            w138=> c0_n77_w138, 
            w139=> c0_n77_w139, 
            w140=> c0_n77_w140, 
            w141=> c0_n77_w141, 
            w142=> c0_n77_w142, 
            w143=> c0_n77_w143, 
            w144=> c0_n77_w144, 
            w145=> c0_n77_w145, 
            w146=> c0_n77_w146, 
            w147=> c0_n77_w147, 
            w148=> c0_n77_w148, 
            w149=> c0_n77_w149, 
            w150=> c0_n77_w150, 
            w151=> c0_n77_w151, 
            w152=> c0_n77_w152, 
            w153=> c0_n77_w153, 
            w154=> c0_n77_w154, 
            w155=> c0_n77_w155, 
            w156=> c0_n77_w156, 
            w157=> c0_n77_w157, 
            w158=> c0_n77_w158, 
            w159=> c0_n77_w159, 
            w160=> c0_n77_w160, 
            w161=> c0_n77_w161, 
            w162=> c0_n77_w162, 
            w163=> c0_n77_w163, 
            w164=> c0_n77_w164, 
            w165=> c0_n77_w165, 
            w166=> c0_n77_w166, 
            w167=> c0_n77_w167, 
            w168=> c0_n77_w168, 
            w169=> c0_n77_w169, 
            w170=> c0_n77_w170, 
            w171=> c0_n77_w171, 
            w172=> c0_n77_w172, 
            w173=> c0_n77_w173, 
            w174=> c0_n77_w174, 
            w175=> c0_n77_w175, 
            w176=> c0_n77_w176, 
            w177=> c0_n77_w177, 
            w178=> c0_n77_w178, 
            w179=> c0_n77_w179, 
            w180=> c0_n77_w180, 
            w181=> c0_n77_w181, 
            w182=> c0_n77_w182, 
            w183=> c0_n77_w183, 
            w184=> c0_n77_w184, 
            w185=> c0_n77_w185, 
            w186=> c0_n77_w186, 
            w187=> c0_n77_w187, 
            w188=> c0_n77_w188, 
            w189=> c0_n77_w189, 
            w190=> c0_n77_w190, 
            w191=> c0_n77_w191, 
            w192=> c0_n77_w192, 
            w193=> c0_n77_w193, 
            w194=> c0_n77_w194, 
            w195=> c0_n77_w195, 
            w196=> c0_n77_w196, 
            w197=> c0_n77_w197, 
            w198=> c0_n77_w198, 
            w199=> c0_n77_w199, 
            w200=> c0_n77_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n77_y
   );           
            
neuron_inst_78: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n78_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n78_w1, 
            w2=> c0_n78_w2, 
            w3=> c0_n78_w3, 
            w4=> c0_n78_w4, 
            w5=> c0_n78_w5, 
            w6=> c0_n78_w6, 
            w7=> c0_n78_w7, 
            w8=> c0_n78_w8, 
            w9=> c0_n78_w9, 
            w10=> c0_n78_w10, 
            w11=> c0_n78_w11, 
            w12=> c0_n78_w12, 
            w13=> c0_n78_w13, 
            w14=> c0_n78_w14, 
            w15=> c0_n78_w15, 
            w16=> c0_n78_w16, 
            w17=> c0_n78_w17, 
            w18=> c0_n78_w18, 
            w19=> c0_n78_w19, 
            w20=> c0_n78_w20, 
            w21=> c0_n78_w21, 
            w22=> c0_n78_w22, 
            w23=> c0_n78_w23, 
            w24=> c0_n78_w24, 
            w25=> c0_n78_w25, 
            w26=> c0_n78_w26, 
            w27=> c0_n78_w27, 
            w28=> c0_n78_w28, 
            w29=> c0_n78_w29, 
            w30=> c0_n78_w30, 
            w31=> c0_n78_w31, 
            w32=> c0_n78_w32, 
            w33=> c0_n78_w33, 
            w34=> c0_n78_w34, 
            w35=> c0_n78_w35, 
            w36=> c0_n78_w36, 
            w37=> c0_n78_w37, 
            w38=> c0_n78_w38, 
            w39=> c0_n78_w39, 
            w40=> c0_n78_w40, 
            w41=> c0_n78_w41, 
            w42=> c0_n78_w42, 
            w43=> c0_n78_w43, 
            w44=> c0_n78_w44, 
            w45=> c0_n78_w45, 
            w46=> c0_n78_w46, 
            w47=> c0_n78_w47, 
            w48=> c0_n78_w48, 
            w49=> c0_n78_w49, 
            w50=> c0_n78_w50, 
            w51=> c0_n78_w51, 
            w52=> c0_n78_w52, 
            w53=> c0_n78_w53, 
            w54=> c0_n78_w54, 
            w55=> c0_n78_w55, 
            w56=> c0_n78_w56, 
            w57=> c0_n78_w57, 
            w58=> c0_n78_w58, 
            w59=> c0_n78_w59, 
            w60=> c0_n78_w60, 
            w61=> c0_n78_w61, 
            w62=> c0_n78_w62, 
            w63=> c0_n78_w63, 
            w64=> c0_n78_w64, 
            w65=> c0_n78_w65, 
            w66=> c0_n78_w66, 
            w67=> c0_n78_w67, 
            w68=> c0_n78_w68, 
            w69=> c0_n78_w69, 
            w70=> c0_n78_w70, 
            w71=> c0_n78_w71, 
            w72=> c0_n78_w72, 
            w73=> c0_n78_w73, 
            w74=> c0_n78_w74, 
            w75=> c0_n78_w75, 
            w76=> c0_n78_w76, 
            w77=> c0_n78_w77, 
            w78=> c0_n78_w78, 
            w79=> c0_n78_w79, 
            w80=> c0_n78_w80, 
            w81=> c0_n78_w81, 
            w82=> c0_n78_w82, 
            w83=> c0_n78_w83, 
            w84=> c0_n78_w84, 
            w85=> c0_n78_w85, 
            w86=> c0_n78_w86, 
            w87=> c0_n78_w87, 
            w88=> c0_n78_w88, 
            w89=> c0_n78_w89, 
            w90=> c0_n78_w90, 
            w91=> c0_n78_w91, 
            w92=> c0_n78_w92, 
            w93=> c0_n78_w93, 
            w94=> c0_n78_w94, 
            w95=> c0_n78_w95, 
            w96=> c0_n78_w96, 
            w97=> c0_n78_w97, 
            w98=> c0_n78_w98, 
            w99=> c0_n78_w99, 
            w100=> c0_n78_w100, 
            w101=> c0_n78_w101, 
            w102=> c0_n78_w102, 
            w103=> c0_n78_w103, 
            w104=> c0_n78_w104, 
            w105=> c0_n78_w105, 
            w106=> c0_n78_w106, 
            w107=> c0_n78_w107, 
            w108=> c0_n78_w108, 
            w109=> c0_n78_w109, 
            w110=> c0_n78_w110, 
            w111=> c0_n78_w111, 
            w112=> c0_n78_w112, 
            w113=> c0_n78_w113, 
            w114=> c0_n78_w114, 
            w115=> c0_n78_w115, 
            w116=> c0_n78_w116, 
            w117=> c0_n78_w117, 
            w118=> c0_n78_w118, 
            w119=> c0_n78_w119, 
            w120=> c0_n78_w120, 
            w121=> c0_n78_w121, 
            w122=> c0_n78_w122, 
            w123=> c0_n78_w123, 
            w124=> c0_n78_w124, 
            w125=> c0_n78_w125, 
            w126=> c0_n78_w126, 
            w127=> c0_n78_w127, 
            w128=> c0_n78_w128, 
            w129=> c0_n78_w129, 
            w130=> c0_n78_w130, 
            w131=> c0_n78_w131, 
            w132=> c0_n78_w132, 
            w133=> c0_n78_w133, 
            w134=> c0_n78_w134, 
            w135=> c0_n78_w135, 
            w136=> c0_n78_w136, 
            w137=> c0_n78_w137, 
            w138=> c0_n78_w138, 
            w139=> c0_n78_w139, 
            w140=> c0_n78_w140, 
            w141=> c0_n78_w141, 
            w142=> c0_n78_w142, 
            w143=> c0_n78_w143, 
            w144=> c0_n78_w144, 
            w145=> c0_n78_w145, 
            w146=> c0_n78_w146, 
            w147=> c0_n78_w147, 
            w148=> c0_n78_w148, 
            w149=> c0_n78_w149, 
            w150=> c0_n78_w150, 
            w151=> c0_n78_w151, 
            w152=> c0_n78_w152, 
            w153=> c0_n78_w153, 
            w154=> c0_n78_w154, 
            w155=> c0_n78_w155, 
            w156=> c0_n78_w156, 
            w157=> c0_n78_w157, 
            w158=> c0_n78_w158, 
            w159=> c0_n78_w159, 
            w160=> c0_n78_w160, 
            w161=> c0_n78_w161, 
            w162=> c0_n78_w162, 
            w163=> c0_n78_w163, 
            w164=> c0_n78_w164, 
            w165=> c0_n78_w165, 
            w166=> c0_n78_w166, 
            w167=> c0_n78_w167, 
            w168=> c0_n78_w168, 
            w169=> c0_n78_w169, 
            w170=> c0_n78_w170, 
            w171=> c0_n78_w171, 
            w172=> c0_n78_w172, 
            w173=> c0_n78_w173, 
            w174=> c0_n78_w174, 
            w175=> c0_n78_w175, 
            w176=> c0_n78_w176, 
            w177=> c0_n78_w177, 
            w178=> c0_n78_w178, 
            w179=> c0_n78_w179, 
            w180=> c0_n78_w180, 
            w181=> c0_n78_w181, 
            w182=> c0_n78_w182, 
            w183=> c0_n78_w183, 
            w184=> c0_n78_w184, 
            w185=> c0_n78_w185, 
            w186=> c0_n78_w186, 
            w187=> c0_n78_w187, 
            w188=> c0_n78_w188, 
            w189=> c0_n78_w189, 
            w190=> c0_n78_w190, 
            w191=> c0_n78_w191, 
            w192=> c0_n78_w192, 
            w193=> c0_n78_w193, 
            w194=> c0_n78_w194, 
            w195=> c0_n78_w195, 
            w196=> c0_n78_w196, 
            w197=> c0_n78_w197, 
            w198=> c0_n78_w198, 
            w199=> c0_n78_w199, 
            w200=> c0_n78_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n78_y
   );           
            
neuron_inst_79: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n79_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n79_w1, 
            w2=> c0_n79_w2, 
            w3=> c0_n79_w3, 
            w4=> c0_n79_w4, 
            w5=> c0_n79_w5, 
            w6=> c0_n79_w6, 
            w7=> c0_n79_w7, 
            w8=> c0_n79_w8, 
            w9=> c0_n79_w9, 
            w10=> c0_n79_w10, 
            w11=> c0_n79_w11, 
            w12=> c0_n79_w12, 
            w13=> c0_n79_w13, 
            w14=> c0_n79_w14, 
            w15=> c0_n79_w15, 
            w16=> c0_n79_w16, 
            w17=> c0_n79_w17, 
            w18=> c0_n79_w18, 
            w19=> c0_n79_w19, 
            w20=> c0_n79_w20, 
            w21=> c0_n79_w21, 
            w22=> c0_n79_w22, 
            w23=> c0_n79_w23, 
            w24=> c0_n79_w24, 
            w25=> c0_n79_w25, 
            w26=> c0_n79_w26, 
            w27=> c0_n79_w27, 
            w28=> c0_n79_w28, 
            w29=> c0_n79_w29, 
            w30=> c0_n79_w30, 
            w31=> c0_n79_w31, 
            w32=> c0_n79_w32, 
            w33=> c0_n79_w33, 
            w34=> c0_n79_w34, 
            w35=> c0_n79_w35, 
            w36=> c0_n79_w36, 
            w37=> c0_n79_w37, 
            w38=> c0_n79_w38, 
            w39=> c0_n79_w39, 
            w40=> c0_n79_w40, 
            w41=> c0_n79_w41, 
            w42=> c0_n79_w42, 
            w43=> c0_n79_w43, 
            w44=> c0_n79_w44, 
            w45=> c0_n79_w45, 
            w46=> c0_n79_w46, 
            w47=> c0_n79_w47, 
            w48=> c0_n79_w48, 
            w49=> c0_n79_w49, 
            w50=> c0_n79_w50, 
            w51=> c0_n79_w51, 
            w52=> c0_n79_w52, 
            w53=> c0_n79_w53, 
            w54=> c0_n79_w54, 
            w55=> c0_n79_w55, 
            w56=> c0_n79_w56, 
            w57=> c0_n79_w57, 
            w58=> c0_n79_w58, 
            w59=> c0_n79_w59, 
            w60=> c0_n79_w60, 
            w61=> c0_n79_w61, 
            w62=> c0_n79_w62, 
            w63=> c0_n79_w63, 
            w64=> c0_n79_w64, 
            w65=> c0_n79_w65, 
            w66=> c0_n79_w66, 
            w67=> c0_n79_w67, 
            w68=> c0_n79_w68, 
            w69=> c0_n79_w69, 
            w70=> c0_n79_w70, 
            w71=> c0_n79_w71, 
            w72=> c0_n79_w72, 
            w73=> c0_n79_w73, 
            w74=> c0_n79_w74, 
            w75=> c0_n79_w75, 
            w76=> c0_n79_w76, 
            w77=> c0_n79_w77, 
            w78=> c0_n79_w78, 
            w79=> c0_n79_w79, 
            w80=> c0_n79_w80, 
            w81=> c0_n79_w81, 
            w82=> c0_n79_w82, 
            w83=> c0_n79_w83, 
            w84=> c0_n79_w84, 
            w85=> c0_n79_w85, 
            w86=> c0_n79_w86, 
            w87=> c0_n79_w87, 
            w88=> c0_n79_w88, 
            w89=> c0_n79_w89, 
            w90=> c0_n79_w90, 
            w91=> c0_n79_w91, 
            w92=> c0_n79_w92, 
            w93=> c0_n79_w93, 
            w94=> c0_n79_w94, 
            w95=> c0_n79_w95, 
            w96=> c0_n79_w96, 
            w97=> c0_n79_w97, 
            w98=> c0_n79_w98, 
            w99=> c0_n79_w99, 
            w100=> c0_n79_w100, 
            w101=> c0_n79_w101, 
            w102=> c0_n79_w102, 
            w103=> c0_n79_w103, 
            w104=> c0_n79_w104, 
            w105=> c0_n79_w105, 
            w106=> c0_n79_w106, 
            w107=> c0_n79_w107, 
            w108=> c0_n79_w108, 
            w109=> c0_n79_w109, 
            w110=> c0_n79_w110, 
            w111=> c0_n79_w111, 
            w112=> c0_n79_w112, 
            w113=> c0_n79_w113, 
            w114=> c0_n79_w114, 
            w115=> c0_n79_w115, 
            w116=> c0_n79_w116, 
            w117=> c0_n79_w117, 
            w118=> c0_n79_w118, 
            w119=> c0_n79_w119, 
            w120=> c0_n79_w120, 
            w121=> c0_n79_w121, 
            w122=> c0_n79_w122, 
            w123=> c0_n79_w123, 
            w124=> c0_n79_w124, 
            w125=> c0_n79_w125, 
            w126=> c0_n79_w126, 
            w127=> c0_n79_w127, 
            w128=> c0_n79_w128, 
            w129=> c0_n79_w129, 
            w130=> c0_n79_w130, 
            w131=> c0_n79_w131, 
            w132=> c0_n79_w132, 
            w133=> c0_n79_w133, 
            w134=> c0_n79_w134, 
            w135=> c0_n79_w135, 
            w136=> c0_n79_w136, 
            w137=> c0_n79_w137, 
            w138=> c0_n79_w138, 
            w139=> c0_n79_w139, 
            w140=> c0_n79_w140, 
            w141=> c0_n79_w141, 
            w142=> c0_n79_w142, 
            w143=> c0_n79_w143, 
            w144=> c0_n79_w144, 
            w145=> c0_n79_w145, 
            w146=> c0_n79_w146, 
            w147=> c0_n79_w147, 
            w148=> c0_n79_w148, 
            w149=> c0_n79_w149, 
            w150=> c0_n79_w150, 
            w151=> c0_n79_w151, 
            w152=> c0_n79_w152, 
            w153=> c0_n79_w153, 
            w154=> c0_n79_w154, 
            w155=> c0_n79_w155, 
            w156=> c0_n79_w156, 
            w157=> c0_n79_w157, 
            w158=> c0_n79_w158, 
            w159=> c0_n79_w159, 
            w160=> c0_n79_w160, 
            w161=> c0_n79_w161, 
            w162=> c0_n79_w162, 
            w163=> c0_n79_w163, 
            w164=> c0_n79_w164, 
            w165=> c0_n79_w165, 
            w166=> c0_n79_w166, 
            w167=> c0_n79_w167, 
            w168=> c0_n79_w168, 
            w169=> c0_n79_w169, 
            w170=> c0_n79_w170, 
            w171=> c0_n79_w171, 
            w172=> c0_n79_w172, 
            w173=> c0_n79_w173, 
            w174=> c0_n79_w174, 
            w175=> c0_n79_w175, 
            w176=> c0_n79_w176, 
            w177=> c0_n79_w177, 
            w178=> c0_n79_w178, 
            w179=> c0_n79_w179, 
            w180=> c0_n79_w180, 
            w181=> c0_n79_w181, 
            w182=> c0_n79_w182, 
            w183=> c0_n79_w183, 
            w184=> c0_n79_w184, 
            w185=> c0_n79_w185, 
            w186=> c0_n79_w186, 
            w187=> c0_n79_w187, 
            w188=> c0_n79_w188, 
            w189=> c0_n79_w189, 
            w190=> c0_n79_w190, 
            w191=> c0_n79_w191, 
            w192=> c0_n79_w192, 
            w193=> c0_n79_w193, 
            w194=> c0_n79_w194, 
            w195=> c0_n79_w195, 
            w196=> c0_n79_w196, 
            w197=> c0_n79_w197, 
            w198=> c0_n79_w198, 
            w199=> c0_n79_w199, 
            w200=> c0_n79_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n79_y
   );           
            
neuron_inst_80: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n80_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n80_w1, 
            w2=> c0_n80_w2, 
            w3=> c0_n80_w3, 
            w4=> c0_n80_w4, 
            w5=> c0_n80_w5, 
            w6=> c0_n80_w6, 
            w7=> c0_n80_w7, 
            w8=> c0_n80_w8, 
            w9=> c0_n80_w9, 
            w10=> c0_n80_w10, 
            w11=> c0_n80_w11, 
            w12=> c0_n80_w12, 
            w13=> c0_n80_w13, 
            w14=> c0_n80_w14, 
            w15=> c0_n80_w15, 
            w16=> c0_n80_w16, 
            w17=> c0_n80_w17, 
            w18=> c0_n80_w18, 
            w19=> c0_n80_w19, 
            w20=> c0_n80_w20, 
            w21=> c0_n80_w21, 
            w22=> c0_n80_w22, 
            w23=> c0_n80_w23, 
            w24=> c0_n80_w24, 
            w25=> c0_n80_w25, 
            w26=> c0_n80_w26, 
            w27=> c0_n80_w27, 
            w28=> c0_n80_w28, 
            w29=> c0_n80_w29, 
            w30=> c0_n80_w30, 
            w31=> c0_n80_w31, 
            w32=> c0_n80_w32, 
            w33=> c0_n80_w33, 
            w34=> c0_n80_w34, 
            w35=> c0_n80_w35, 
            w36=> c0_n80_w36, 
            w37=> c0_n80_w37, 
            w38=> c0_n80_w38, 
            w39=> c0_n80_w39, 
            w40=> c0_n80_w40, 
            w41=> c0_n80_w41, 
            w42=> c0_n80_w42, 
            w43=> c0_n80_w43, 
            w44=> c0_n80_w44, 
            w45=> c0_n80_w45, 
            w46=> c0_n80_w46, 
            w47=> c0_n80_w47, 
            w48=> c0_n80_w48, 
            w49=> c0_n80_w49, 
            w50=> c0_n80_w50, 
            w51=> c0_n80_w51, 
            w52=> c0_n80_w52, 
            w53=> c0_n80_w53, 
            w54=> c0_n80_w54, 
            w55=> c0_n80_w55, 
            w56=> c0_n80_w56, 
            w57=> c0_n80_w57, 
            w58=> c0_n80_w58, 
            w59=> c0_n80_w59, 
            w60=> c0_n80_w60, 
            w61=> c0_n80_w61, 
            w62=> c0_n80_w62, 
            w63=> c0_n80_w63, 
            w64=> c0_n80_w64, 
            w65=> c0_n80_w65, 
            w66=> c0_n80_w66, 
            w67=> c0_n80_w67, 
            w68=> c0_n80_w68, 
            w69=> c0_n80_w69, 
            w70=> c0_n80_w70, 
            w71=> c0_n80_w71, 
            w72=> c0_n80_w72, 
            w73=> c0_n80_w73, 
            w74=> c0_n80_w74, 
            w75=> c0_n80_w75, 
            w76=> c0_n80_w76, 
            w77=> c0_n80_w77, 
            w78=> c0_n80_w78, 
            w79=> c0_n80_w79, 
            w80=> c0_n80_w80, 
            w81=> c0_n80_w81, 
            w82=> c0_n80_w82, 
            w83=> c0_n80_w83, 
            w84=> c0_n80_w84, 
            w85=> c0_n80_w85, 
            w86=> c0_n80_w86, 
            w87=> c0_n80_w87, 
            w88=> c0_n80_w88, 
            w89=> c0_n80_w89, 
            w90=> c0_n80_w90, 
            w91=> c0_n80_w91, 
            w92=> c0_n80_w92, 
            w93=> c0_n80_w93, 
            w94=> c0_n80_w94, 
            w95=> c0_n80_w95, 
            w96=> c0_n80_w96, 
            w97=> c0_n80_w97, 
            w98=> c0_n80_w98, 
            w99=> c0_n80_w99, 
            w100=> c0_n80_w100, 
            w101=> c0_n80_w101, 
            w102=> c0_n80_w102, 
            w103=> c0_n80_w103, 
            w104=> c0_n80_w104, 
            w105=> c0_n80_w105, 
            w106=> c0_n80_w106, 
            w107=> c0_n80_w107, 
            w108=> c0_n80_w108, 
            w109=> c0_n80_w109, 
            w110=> c0_n80_w110, 
            w111=> c0_n80_w111, 
            w112=> c0_n80_w112, 
            w113=> c0_n80_w113, 
            w114=> c0_n80_w114, 
            w115=> c0_n80_w115, 
            w116=> c0_n80_w116, 
            w117=> c0_n80_w117, 
            w118=> c0_n80_w118, 
            w119=> c0_n80_w119, 
            w120=> c0_n80_w120, 
            w121=> c0_n80_w121, 
            w122=> c0_n80_w122, 
            w123=> c0_n80_w123, 
            w124=> c0_n80_w124, 
            w125=> c0_n80_w125, 
            w126=> c0_n80_w126, 
            w127=> c0_n80_w127, 
            w128=> c0_n80_w128, 
            w129=> c0_n80_w129, 
            w130=> c0_n80_w130, 
            w131=> c0_n80_w131, 
            w132=> c0_n80_w132, 
            w133=> c0_n80_w133, 
            w134=> c0_n80_w134, 
            w135=> c0_n80_w135, 
            w136=> c0_n80_w136, 
            w137=> c0_n80_w137, 
            w138=> c0_n80_w138, 
            w139=> c0_n80_w139, 
            w140=> c0_n80_w140, 
            w141=> c0_n80_w141, 
            w142=> c0_n80_w142, 
            w143=> c0_n80_w143, 
            w144=> c0_n80_w144, 
            w145=> c0_n80_w145, 
            w146=> c0_n80_w146, 
            w147=> c0_n80_w147, 
            w148=> c0_n80_w148, 
            w149=> c0_n80_w149, 
            w150=> c0_n80_w150, 
            w151=> c0_n80_w151, 
            w152=> c0_n80_w152, 
            w153=> c0_n80_w153, 
            w154=> c0_n80_w154, 
            w155=> c0_n80_w155, 
            w156=> c0_n80_w156, 
            w157=> c0_n80_w157, 
            w158=> c0_n80_w158, 
            w159=> c0_n80_w159, 
            w160=> c0_n80_w160, 
            w161=> c0_n80_w161, 
            w162=> c0_n80_w162, 
            w163=> c0_n80_w163, 
            w164=> c0_n80_w164, 
            w165=> c0_n80_w165, 
            w166=> c0_n80_w166, 
            w167=> c0_n80_w167, 
            w168=> c0_n80_w168, 
            w169=> c0_n80_w169, 
            w170=> c0_n80_w170, 
            w171=> c0_n80_w171, 
            w172=> c0_n80_w172, 
            w173=> c0_n80_w173, 
            w174=> c0_n80_w174, 
            w175=> c0_n80_w175, 
            w176=> c0_n80_w176, 
            w177=> c0_n80_w177, 
            w178=> c0_n80_w178, 
            w179=> c0_n80_w179, 
            w180=> c0_n80_w180, 
            w181=> c0_n80_w181, 
            w182=> c0_n80_w182, 
            w183=> c0_n80_w183, 
            w184=> c0_n80_w184, 
            w185=> c0_n80_w185, 
            w186=> c0_n80_w186, 
            w187=> c0_n80_w187, 
            w188=> c0_n80_w188, 
            w189=> c0_n80_w189, 
            w190=> c0_n80_w190, 
            w191=> c0_n80_w191, 
            w192=> c0_n80_w192, 
            w193=> c0_n80_w193, 
            w194=> c0_n80_w194, 
            w195=> c0_n80_w195, 
            w196=> c0_n80_w196, 
            w197=> c0_n80_w197, 
            w198=> c0_n80_w198, 
            w199=> c0_n80_w199, 
            w200=> c0_n80_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n80_y
   );           
            
neuron_inst_81: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n81_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n81_w1, 
            w2=> c0_n81_w2, 
            w3=> c0_n81_w3, 
            w4=> c0_n81_w4, 
            w5=> c0_n81_w5, 
            w6=> c0_n81_w6, 
            w7=> c0_n81_w7, 
            w8=> c0_n81_w8, 
            w9=> c0_n81_w9, 
            w10=> c0_n81_w10, 
            w11=> c0_n81_w11, 
            w12=> c0_n81_w12, 
            w13=> c0_n81_w13, 
            w14=> c0_n81_w14, 
            w15=> c0_n81_w15, 
            w16=> c0_n81_w16, 
            w17=> c0_n81_w17, 
            w18=> c0_n81_w18, 
            w19=> c0_n81_w19, 
            w20=> c0_n81_w20, 
            w21=> c0_n81_w21, 
            w22=> c0_n81_w22, 
            w23=> c0_n81_w23, 
            w24=> c0_n81_w24, 
            w25=> c0_n81_w25, 
            w26=> c0_n81_w26, 
            w27=> c0_n81_w27, 
            w28=> c0_n81_w28, 
            w29=> c0_n81_w29, 
            w30=> c0_n81_w30, 
            w31=> c0_n81_w31, 
            w32=> c0_n81_w32, 
            w33=> c0_n81_w33, 
            w34=> c0_n81_w34, 
            w35=> c0_n81_w35, 
            w36=> c0_n81_w36, 
            w37=> c0_n81_w37, 
            w38=> c0_n81_w38, 
            w39=> c0_n81_w39, 
            w40=> c0_n81_w40, 
            w41=> c0_n81_w41, 
            w42=> c0_n81_w42, 
            w43=> c0_n81_w43, 
            w44=> c0_n81_w44, 
            w45=> c0_n81_w45, 
            w46=> c0_n81_w46, 
            w47=> c0_n81_w47, 
            w48=> c0_n81_w48, 
            w49=> c0_n81_w49, 
            w50=> c0_n81_w50, 
            w51=> c0_n81_w51, 
            w52=> c0_n81_w52, 
            w53=> c0_n81_w53, 
            w54=> c0_n81_w54, 
            w55=> c0_n81_w55, 
            w56=> c0_n81_w56, 
            w57=> c0_n81_w57, 
            w58=> c0_n81_w58, 
            w59=> c0_n81_w59, 
            w60=> c0_n81_w60, 
            w61=> c0_n81_w61, 
            w62=> c0_n81_w62, 
            w63=> c0_n81_w63, 
            w64=> c0_n81_w64, 
            w65=> c0_n81_w65, 
            w66=> c0_n81_w66, 
            w67=> c0_n81_w67, 
            w68=> c0_n81_w68, 
            w69=> c0_n81_w69, 
            w70=> c0_n81_w70, 
            w71=> c0_n81_w71, 
            w72=> c0_n81_w72, 
            w73=> c0_n81_w73, 
            w74=> c0_n81_w74, 
            w75=> c0_n81_w75, 
            w76=> c0_n81_w76, 
            w77=> c0_n81_w77, 
            w78=> c0_n81_w78, 
            w79=> c0_n81_w79, 
            w80=> c0_n81_w80, 
            w81=> c0_n81_w81, 
            w82=> c0_n81_w82, 
            w83=> c0_n81_w83, 
            w84=> c0_n81_w84, 
            w85=> c0_n81_w85, 
            w86=> c0_n81_w86, 
            w87=> c0_n81_w87, 
            w88=> c0_n81_w88, 
            w89=> c0_n81_w89, 
            w90=> c0_n81_w90, 
            w91=> c0_n81_w91, 
            w92=> c0_n81_w92, 
            w93=> c0_n81_w93, 
            w94=> c0_n81_w94, 
            w95=> c0_n81_w95, 
            w96=> c0_n81_w96, 
            w97=> c0_n81_w97, 
            w98=> c0_n81_w98, 
            w99=> c0_n81_w99, 
            w100=> c0_n81_w100, 
            w101=> c0_n81_w101, 
            w102=> c0_n81_w102, 
            w103=> c0_n81_w103, 
            w104=> c0_n81_w104, 
            w105=> c0_n81_w105, 
            w106=> c0_n81_w106, 
            w107=> c0_n81_w107, 
            w108=> c0_n81_w108, 
            w109=> c0_n81_w109, 
            w110=> c0_n81_w110, 
            w111=> c0_n81_w111, 
            w112=> c0_n81_w112, 
            w113=> c0_n81_w113, 
            w114=> c0_n81_w114, 
            w115=> c0_n81_w115, 
            w116=> c0_n81_w116, 
            w117=> c0_n81_w117, 
            w118=> c0_n81_w118, 
            w119=> c0_n81_w119, 
            w120=> c0_n81_w120, 
            w121=> c0_n81_w121, 
            w122=> c0_n81_w122, 
            w123=> c0_n81_w123, 
            w124=> c0_n81_w124, 
            w125=> c0_n81_w125, 
            w126=> c0_n81_w126, 
            w127=> c0_n81_w127, 
            w128=> c0_n81_w128, 
            w129=> c0_n81_w129, 
            w130=> c0_n81_w130, 
            w131=> c0_n81_w131, 
            w132=> c0_n81_w132, 
            w133=> c0_n81_w133, 
            w134=> c0_n81_w134, 
            w135=> c0_n81_w135, 
            w136=> c0_n81_w136, 
            w137=> c0_n81_w137, 
            w138=> c0_n81_w138, 
            w139=> c0_n81_w139, 
            w140=> c0_n81_w140, 
            w141=> c0_n81_w141, 
            w142=> c0_n81_w142, 
            w143=> c0_n81_w143, 
            w144=> c0_n81_w144, 
            w145=> c0_n81_w145, 
            w146=> c0_n81_w146, 
            w147=> c0_n81_w147, 
            w148=> c0_n81_w148, 
            w149=> c0_n81_w149, 
            w150=> c0_n81_w150, 
            w151=> c0_n81_w151, 
            w152=> c0_n81_w152, 
            w153=> c0_n81_w153, 
            w154=> c0_n81_w154, 
            w155=> c0_n81_w155, 
            w156=> c0_n81_w156, 
            w157=> c0_n81_w157, 
            w158=> c0_n81_w158, 
            w159=> c0_n81_w159, 
            w160=> c0_n81_w160, 
            w161=> c0_n81_w161, 
            w162=> c0_n81_w162, 
            w163=> c0_n81_w163, 
            w164=> c0_n81_w164, 
            w165=> c0_n81_w165, 
            w166=> c0_n81_w166, 
            w167=> c0_n81_w167, 
            w168=> c0_n81_w168, 
            w169=> c0_n81_w169, 
            w170=> c0_n81_w170, 
            w171=> c0_n81_w171, 
            w172=> c0_n81_w172, 
            w173=> c0_n81_w173, 
            w174=> c0_n81_w174, 
            w175=> c0_n81_w175, 
            w176=> c0_n81_w176, 
            w177=> c0_n81_w177, 
            w178=> c0_n81_w178, 
            w179=> c0_n81_w179, 
            w180=> c0_n81_w180, 
            w181=> c0_n81_w181, 
            w182=> c0_n81_w182, 
            w183=> c0_n81_w183, 
            w184=> c0_n81_w184, 
            w185=> c0_n81_w185, 
            w186=> c0_n81_w186, 
            w187=> c0_n81_w187, 
            w188=> c0_n81_w188, 
            w189=> c0_n81_w189, 
            w190=> c0_n81_w190, 
            w191=> c0_n81_w191, 
            w192=> c0_n81_w192, 
            w193=> c0_n81_w193, 
            w194=> c0_n81_w194, 
            w195=> c0_n81_w195, 
            w196=> c0_n81_w196, 
            w197=> c0_n81_w197, 
            w198=> c0_n81_w198, 
            w199=> c0_n81_w199, 
            w200=> c0_n81_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n81_y
   );           
            
neuron_inst_82: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n82_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n82_w1, 
            w2=> c0_n82_w2, 
            w3=> c0_n82_w3, 
            w4=> c0_n82_w4, 
            w5=> c0_n82_w5, 
            w6=> c0_n82_w6, 
            w7=> c0_n82_w7, 
            w8=> c0_n82_w8, 
            w9=> c0_n82_w9, 
            w10=> c0_n82_w10, 
            w11=> c0_n82_w11, 
            w12=> c0_n82_w12, 
            w13=> c0_n82_w13, 
            w14=> c0_n82_w14, 
            w15=> c0_n82_w15, 
            w16=> c0_n82_w16, 
            w17=> c0_n82_w17, 
            w18=> c0_n82_w18, 
            w19=> c0_n82_w19, 
            w20=> c0_n82_w20, 
            w21=> c0_n82_w21, 
            w22=> c0_n82_w22, 
            w23=> c0_n82_w23, 
            w24=> c0_n82_w24, 
            w25=> c0_n82_w25, 
            w26=> c0_n82_w26, 
            w27=> c0_n82_w27, 
            w28=> c0_n82_w28, 
            w29=> c0_n82_w29, 
            w30=> c0_n82_w30, 
            w31=> c0_n82_w31, 
            w32=> c0_n82_w32, 
            w33=> c0_n82_w33, 
            w34=> c0_n82_w34, 
            w35=> c0_n82_w35, 
            w36=> c0_n82_w36, 
            w37=> c0_n82_w37, 
            w38=> c0_n82_w38, 
            w39=> c0_n82_w39, 
            w40=> c0_n82_w40, 
            w41=> c0_n82_w41, 
            w42=> c0_n82_w42, 
            w43=> c0_n82_w43, 
            w44=> c0_n82_w44, 
            w45=> c0_n82_w45, 
            w46=> c0_n82_w46, 
            w47=> c0_n82_w47, 
            w48=> c0_n82_w48, 
            w49=> c0_n82_w49, 
            w50=> c0_n82_w50, 
            w51=> c0_n82_w51, 
            w52=> c0_n82_w52, 
            w53=> c0_n82_w53, 
            w54=> c0_n82_w54, 
            w55=> c0_n82_w55, 
            w56=> c0_n82_w56, 
            w57=> c0_n82_w57, 
            w58=> c0_n82_w58, 
            w59=> c0_n82_w59, 
            w60=> c0_n82_w60, 
            w61=> c0_n82_w61, 
            w62=> c0_n82_w62, 
            w63=> c0_n82_w63, 
            w64=> c0_n82_w64, 
            w65=> c0_n82_w65, 
            w66=> c0_n82_w66, 
            w67=> c0_n82_w67, 
            w68=> c0_n82_w68, 
            w69=> c0_n82_w69, 
            w70=> c0_n82_w70, 
            w71=> c0_n82_w71, 
            w72=> c0_n82_w72, 
            w73=> c0_n82_w73, 
            w74=> c0_n82_w74, 
            w75=> c0_n82_w75, 
            w76=> c0_n82_w76, 
            w77=> c0_n82_w77, 
            w78=> c0_n82_w78, 
            w79=> c0_n82_w79, 
            w80=> c0_n82_w80, 
            w81=> c0_n82_w81, 
            w82=> c0_n82_w82, 
            w83=> c0_n82_w83, 
            w84=> c0_n82_w84, 
            w85=> c0_n82_w85, 
            w86=> c0_n82_w86, 
            w87=> c0_n82_w87, 
            w88=> c0_n82_w88, 
            w89=> c0_n82_w89, 
            w90=> c0_n82_w90, 
            w91=> c0_n82_w91, 
            w92=> c0_n82_w92, 
            w93=> c0_n82_w93, 
            w94=> c0_n82_w94, 
            w95=> c0_n82_w95, 
            w96=> c0_n82_w96, 
            w97=> c0_n82_w97, 
            w98=> c0_n82_w98, 
            w99=> c0_n82_w99, 
            w100=> c0_n82_w100, 
            w101=> c0_n82_w101, 
            w102=> c0_n82_w102, 
            w103=> c0_n82_w103, 
            w104=> c0_n82_w104, 
            w105=> c0_n82_w105, 
            w106=> c0_n82_w106, 
            w107=> c0_n82_w107, 
            w108=> c0_n82_w108, 
            w109=> c0_n82_w109, 
            w110=> c0_n82_w110, 
            w111=> c0_n82_w111, 
            w112=> c0_n82_w112, 
            w113=> c0_n82_w113, 
            w114=> c0_n82_w114, 
            w115=> c0_n82_w115, 
            w116=> c0_n82_w116, 
            w117=> c0_n82_w117, 
            w118=> c0_n82_w118, 
            w119=> c0_n82_w119, 
            w120=> c0_n82_w120, 
            w121=> c0_n82_w121, 
            w122=> c0_n82_w122, 
            w123=> c0_n82_w123, 
            w124=> c0_n82_w124, 
            w125=> c0_n82_w125, 
            w126=> c0_n82_w126, 
            w127=> c0_n82_w127, 
            w128=> c0_n82_w128, 
            w129=> c0_n82_w129, 
            w130=> c0_n82_w130, 
            w131=> c0_n82_w131, 
            w132=> c0_n82_w132, 
            w133=> c0_n82_w133, 
            w134=> c0_n82_w134, 
            w135=> c0_n82_w135, 
            w136=> c0_n82_w136, 
            w137=> c0_n82_w137, 
            w138=> c0_n82_w138, 
            w139=> c0_n82_w139, 
            w140=> c0_n82_w140, 
            w141=> c0_n82_w141, 
            w142=> c0_n82_w142, 
            w143=> c0_n82_w143, 
            w144=> c0_n82_w144, 
            w145=> c0_n82_w145, 
            w146=> c0_n82_w146, 
            w147=> c0_n82_w147, 
            w148=> c0_n82_w148, 
            w149=> c0_n82_w149, 
            w150=> c0_n82_w150, 
            w151=> c0_n82_w151, 
            w152=> c0_n82_w152, 
            w153=> c0_n82_w153, 
            w154=> c0_n82_w154, 
            w155=> c0_n82_w155, 
            w156=> c0_n82_w156, 
            w157=> c0_n82_w157, 
            w158=> c0_n82_w158, 
            w159=> c0_n82_w159, 
            w160=> c0_n82_w160, 
            w161=> c0_n82_w161, 
            w162=> c0_n82_w162, 
            w163=> c0_n82_w163, 
            w164=> c0_n82_w164, 
            w165=> c0_n82_w165, 
            w166=> c0_n82_w166, 
            w167=> c0_n82_w167, 
            w168=> c0_n82_w168, 
            w169=> c0_n82_w169, 
            w170=> c0_n82_w170, 
            w171=> c0_n82_w171, 
            w172=> c0_n82_w172, 
            w173=> c0_n82_w173, 
            w174=> c0_n82_w174, 
            w175=> c0_n82_w175, 
            w176=> c0_n82_w176, 
            w177=> c0_n82_w177, 
            w178=> c0_n82_w178, 
            w179=> c0_n82_w179, 
            w180=> c0_n82_w180, 
            w181=> c0_n82_w181, 
            w182=> c0_n82_w182, 
            w183=> c0_n82_w183, 
            w184=> c0_n82_w184, 
            w185=> c0_n82_w185, 
            w186=> c0_n82_w186, 
            w187=> c0_n82_w187, 
            w188=> c0_n82_w188, 
            w189=> c0_n82_w189, 
            w190=> c0_n82_w190, 
            w191=> c0_n82_w191, 
            w192=> c0_n82_w192, 
            w193=> c0_n82_w193, 
            w194=> c0_n82_w194, 
            w195=> c0_n82_w195, 
            w196=> c0_n82_w196, 
            w197=> c0_n82_w197, 
            w198=> c0_n82_w198, 
            w199=> c0_n82_w199, 
            w200=> c0_n82_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n82_y
   );           
            
neuron_inst_83: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n83_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n83_w1, 
            w2=> c0_n83_w2, 
            w3=> c0_n83_w3, 
            w4=> c0_n83_w4, 
            w5=> c0_n83_w5, 
            w6=> c0_n83_w6, 
            w7=> c0_n83_w7, 
            w8=> c0_n83_w8, 
            w9=> c0_n83_w9, 
            w10=> c0_n83_w10, 
            w11=> c0_n83_w11, 
            w12=> c0_n83_w12, 
            w13=> c0_n83_w13, 
            w14=> c0_n83_w14, 
            w15=> c0_n83_w15, 
            w16=> c0_n83_w16, 
            w17=> c0_n83_w17, 
            w18=> c0_n83_w18, 
            w19=> c0_n83_w19, 
            w20=> c0_n83_w20, 
            w21=> c0_n83_w21, 
            w22=> c0_n83_w22, 
            w23=> c0_n83_w23, 
            w24=> c0_n83_w24, 
            w25=> c0_n83_w25, 
            w26=> c0_n83_w26, 
            w27=> c0_n83_w27, 
            w28=> c0_n83_w28, 
            w29=> c0_n83_w29, 
            w30=> c0_n83_w30, 
            w31=> c0_n83_w31, 
            w32=> c0_n83_w32, 
            w33=> c0_n83_w33, 
            w34=> c0_n83_w34, 
            w35=> c0_n83_w35, 
            w36=> c0_n83_w36, 
            w37=> c0_n83_w37, 
            w38=> c0_n83_w38, 
            w39=> c0_n83_w39, 
            w40=> c0_n83_w40, 
            w41=> c0_n83_w41, 
            w42=> c0_n83_w42, 
            w43=> c0_n83_w43, 
            w44=> c0_n83_w44, 
            w45=> c0_n83_w45, 
            w46=> c0_n83_w46, 
            w47=> c0_n83_w47, 
            w48=> c0_n83_w48, 
            w49=> c0_n83_w49, 
            w50=> c0_n83_w50, 
            w51=> c0_n83_w51, 
            w52=> c0_n83_w52, 
            w53=> c0_n83_w53, 
            w54=> c0_n83_w54, 
            w55=> c0_n83_w55, 
            w56=> c0_n83_w56, 
            w57=> c0_n83_w57, 
            w58=> c0_n83_w58, 
            w59=> c0_n83_w59, 
            w60=> c0_n83_w60, 
            w61=> c0_n83_w61, 
            w62=> c0_n83_w62, 
            w63=> c0_n83_w63, 
            w64=> c0_n83_w64, 
            w65=> c0_n83_w65, 
            w66=> c0_n83_w66, 
            w67=> c0_n83_w67, 
            w68=> c0_n83_w68, 
            w69=> c0_n83_w69, 
            w70=> c0_n83_w70, 
            w71=> c0_n83_w71, 
            w72=> c0_n83_w72, 
            w73=> c0_n83_w73, 
            w74=> c0_n83_w74, 
            w75=> c0_n83_w75, 
            w76=> c0_n83_w76, 
            w77=> c0_n83_w77, 
            w78=> c0_n83_w78, 
            w79=> c0_n83_w79, 
            w80=> c0_n83_w80, 
            w81=> c0_n83_w81, 
            w82=> c0_n83_w82, 
            w83=> c0_n83_w83, 
            w84=> c0_n83_w84, 
            w85=> c0_n83_w85, 
            w86=> c0_n83_w86, 
            w87=> c0_n83_w87, 
            w88=> c0_n83_w88, 
            w89=> c0_n83_w89, 
            w90=> c0_n83_w90, 
            w91=> c0_n83_w91, 
            w92=> c0_n83_w92, 
            w93=> c0_n83_w93, 
            w94=> c0_n83_w94, 
            w95=> c0_n83_w95, 
            w96=> c0_n83_w96, 
            w97=> c0_n83_w97, 
            w98=> c0_n83_w98, 
            w99=> c0_n83_w99, 
            w100=> c0_n83_w100, 
            w101=> c0_n83_w101, 
            w102=> c0_n83_w102, 
            w103=> c0_n83_w103, 
            w104=> c0_n83_w104, 
            w105=> c0_n83_w105, 
            w106=> c0_n83_w106, 
            w107=> c0_n83_w107, 
            w108=> c0_n83_w108, 
            w109=> c0_n83_w109, 
            w110=> c0_n83_w110, 
            w111=> c0_n83_w111, 
            w112=> c0_n83_w112, 
            w113=> c0_n83_w113, 
            w114=> c0_n83_w114, 
            w115=> c0_n83_w115, 
            w116=> c0_n83_w116, 
            w117=> c0_n83_w117, 
            w118=> c0_n83_w118, 
            w119=> c0_n83_w119, 
            w120=> c0_n83_w120, 
            w121=> c0_n83_w121, 
            w122=> c0_n83_w122, 
            w123=> c0_n83_w123, 
            w124=> c0_n83_w124, 
            w125=> c0_n83_w125, 
            w126=> c0_n83_w126, 
            w127=> c0_n83_w127, 
            w128=> c0_n83_w128, 
            w129=> c0_n83_w129, 
            w130=> c0_n83_w130, 
            w131=> c0_n83_w131, 
            w132=> c0_n83_w132, 
            w133=> c0_n83_w133, 
            w134=> c0_n83_w134, 
            w135=> c0_n83_w135, 
            w136=> c0_n83_w136, 
            w137=> c0_n83_w137, 
            w138=> c0_n83_w138, 
            w139=> c0_n83_w139, 
            w140=> c0_n83_w140, 
            w141=> c0_n83_w141, 
            w142=> c0_n83_w142, 
            w143=> c0_n83_w143, 
            w144=> c0_n83_w144, 
            w145=> c0_n83_w145, 
            w146=> c0_n83_w146, 
            w147=> c0_n83_w147, 
            w148=> c0_n83_w148, 
            w149=> c0_n83_w149, 
            w150=> c0_n83_w150, 
            w151=> c0_n83_w151, 
            w152=> c0_n83_w152, 
            w153=> c0_n83_w153, 
            w154=> c0_n83_w154, 
            w155=> c0_n83_w155, 
            w156=> c0_n83_w156, 
            w157=> c0_n83_w157, 
            w158=> c0_n83_w158, 
            w159=> c0_n83_w159, 
            w160=> c0_n83_w160, 
            w161=> c0_n83_w161, 
            w162=> c0_n83_w162, 
            w163=> c0_n83_w163, 
            w164=> c0_n83_w164, 
            w165=> c0_n83_w165, 
            w166=> c0_n83_w166, 
            w167=> c0_n83_w167, 
            w168=> c0_n83_w168, 
            w169=> c0_n83_w169, 
            w170=> c0_n83_w170, 
            w171=> c0_n83_w171, 
            w172=> c0_n83_w172, 
            w173=> c0_n83_w173, 
            w174=> c0_n83_w174, 
            w175=> c0_n83_w175, 
            w176=> c0_n83_w176, 
            w177=> c0_n83_w177, 
            w178=> c0_n83_w178, 
            w179=> c0_n83_w179, 
            w180=> c0_n83_w180, 
            w181=> c0_n83_w181, 
            w182=> c0_n83_w182, 
            w183=> c0_n83_w183, 
            w184=> c0_n83_w184, 
            w185=> c0_n83_w185, 
            w186=> c0_n83_w186, 
            w187=> c0_n83_w187, 
            w188=> c0_n83_w188, 
            w189=> c0_n83_w189, 
            w190=> c0_n83_w190, 
            w191=> c0_n83_w191, 
            w192=> c0_n83_w192, 
            w193=> c0_n83_w193, 
            w194=> c0_n83_w194, 
            w195=> c0_n83_w195, 
            w196=> c0_n83_w196, 
            w197=> c0_n83_w197, 
            w198=> c0_n83_w198, 
            w199=> c0_n83_w199, 
            w200=> c0_n83_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n83_y
   );           
            
neuron_inst_84: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n84_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n84_w1, 
            w2=> c0_n84_w2, 
            w3=> c0_n84_w3, 
            w4=> c0_n84_w4, 
            w5=> c0_n84_w5, 
            w6=> c0_n84_w6, 
            w7=> c0_n84_w7, 
            w8=> c0_n84_w8, 
            w9=> c0_n84_w9, 
            w10=> c0_n84_w10, 
            w11=> c0_n84_w11, 
            w12=> c0_n84_w12, 
            w13=> c0_n84_w13, 
            w14=> c0_n84_w14, 
            w15=> c0_n84_w15, 
            w16=> c0_n84_w16, 
            w17=> c0_n84_w17, 
            w18=> c0_n84_w18, 
            w19=> c0_n84_w19, 
            w20=> c0_n84_w20, 
            w21=> c0_n84_w21, 
            w22=> c0_n84_w22, 
            w23=> c0_n84_w23, 
            w24=> c0_n84_w24, 
            w25=> c0_n84_w25, 
            w26=> c0_n84_w26, 
            w27=> c0_n84_w27, 
            w28=> c0_n84_w28, 
            w29=> c0_n84_w29, 
            w30=> c0_n84_w30, 
            w31=> c0_n84_w31, 
            w32=> c0_n84_w32, 
            w33=> c0_n84_w33, 
            w34=> c0_n84_w34, 
            w35=> c0_n84_w35, 
            w36=> c0_n84_w36, 
            w37=> c0_n84_w37, 
            w38=> c0_n84_w38, 
            w39=> c0_n84_w39, 
            w40=> c0_n84_w40, 
            w41=> c0_n84_w41, 
            w42=> c0_n84_w42, 
            w43=> c0_n84_w43, 
            w44=> c0_n84_w44, 
            w45=> c0_n84_w45, 
            w46=> c0_n84_w46, 
            w47=> c0_n84_w47, 
            w48=> c0_n84_w48, 
            w49=> c0_n84_w49, 
            w50=> c0_n84_w50, 
            w51=> c0_n84_w51, 
            w52=> c0_n84_w52, 
            w53=> c0_n84_w53, 
            w54=> c0_n84_w54, 
            w55=> c0_n84_w55, 
            w56=> c0_n84_w56, 
            w57=> c0_n84_w57, 
            w58=> c0_n84_w58, 
            w59=> c0_n84_w59, 
            w60=> c0_n84_w60, 
            w61=> c0_n84_w61, 
            w62=> c0_n84_w62, 
            w63=> c0_n84_w63, 
            w64=> c0_n84_w64, 
            w65=> c0_n84_w65, 
            w66=> c0_n84_w66, 
            w67=> c0_n84_w67, 
            w68=> c0_n84_w68, 
            w69=> c0_n84_w69, 
            w70=> c0_n84_w70, 
            w71=> c0_n84_w71, 
            w72=> c0_n84_w72, 
            w73=> c0_n84_w73, 
            w74=> c0_n84_w74, 
            w75=> c0_n84_w75, 
            w76=> c0_n84_w76, 
            w77=> c0_n84_w77, 
            w78=> c0_n84_w78, 
            w79=> c0_n84_w79, 
            w80=> c0_n84_w80, 
            w81=> c0_n84_w81, 
            w82=> c0_n84_w82, 
            w83=> c0_n84_w83, 
            w84=> c0_n84_w84, 
            w85=> c0_n84_w85, 
            w86=> c0_n84_w86, 
            w87=> c0_n84_w87, 
            w88=> c0_n84_w88, 
            w89=> c0_n84_w89, 
            w90=> c0_n84_w90, 
            w91=> c0_n84_w91, 
            w92=> c0_n84_w92, 
            w93=> c0_n84_w93, 
            w94=> c0_n84_w94, 
            w95=> c0_n84_w95, 
            w96=> c0_n84_w96, 
            w97=> c0_n84_w97, 
            w98=> c0_n84_w98, 
            w99=> c0_n84_w99, 
            w100=> c0_n84_w100, 
            w101=> c0_n84_w101, 
            w102=> c0_n84_w102, 
            w103=> c0_n84_w103, 
            w104=> c0_n84_w104, 
            w105=> c0_n84_w105, 
            w106=> c0_n84_w106, 
            w107=> c0_n84_w107, 
            w108=> c0_n84_w108, 
            w109=> c0_n84_w109, 
            w110=> c0_n84_w110, 
            w111=> c0_n84_w111, 
            w112=> c0_n84_w112, 
            w113=> c0_n84_w113, 
            w114=> c0_n84_w114, 
            w115=> c0_n84_w115, 
            w116=> c0_n84_w116, 
            w117=> c0_n84_w117, 
            w118=> c0_n84_w118, 
            w119=> c0_n84_w119, 
            w120=> c0_n84_w120, 
            w121=> c0_n84_w121, 
            w122=> c0_n84_w122, 
            w123=> c0_n84_w123, 
            w124=> c0_n84_w124, 
            w125=> c0_n84_w125, 
            w126=> c0_n84_w126, 
            w127=> c0_n84_w127, 
            w128=> c0_n84_w128, 
            w129=> c0_n84_w129, 
            w130=> c0_n84_w130, 
            w131=> c0_n84_w131, 
            w132=> c0_n84_w132, 
            w133=> c0_n84_w133, 
            w134=> c0_n84_w134, 
            w135=> c0_n84_w135, 
            w136=> c0_n84_w136, 
            w137=> c0_n84_w137, 
            w138=> c0_n84_w138, 
            w139=> c0_n84_w139, 
            w140=> c0_n84_w140, 
            w141=> c0_n84_w141, 
            w142=> c0_n84_w142, 
            w143=> c0_n84_w143, 
            w144=> c0_n84_w144, 
            w145=> c0_n84_w145, 
            w146=> c0_n84_w146, 
            w147=> c0_n84_w147, 
            w148=> c0_n84_w148, 
            w149=> c0_n84_w149, 
            w150=> c0_n84_w150, 
            w151=> c0_n84_w151, 
            w152=> c0_n84_w152, 
            w153=> c0_n84_w153, 
            w154=> c0_n84_w154, 
            w155=> c0_n84_w155, 
            w156=> c0_n84_w156, 
            w157=> c0_n84_w157, 
            w158=> c0_n84_w158, 
            w159=> c0_n84_w159, 
            w160=> c0_n84_w160, 
            w161=> c0_n84_w161, 
            w162=> c0_n84_w162, 
            w163=> c0_n84_w163, 
            w164=> c0_n84_w164, 
            w165=> c0_n84_w165, 
            w166=> c0_n84_w166, 
            w167=> c0_n84_w167, 
            w168=> c0_n84_w168, 
            w169=> c0_n84_w169, 
            w170=> c0_n84_w170, 
            w171=> c0_n84_w171, 
            w172=> c0_n84_w172, 
            w173=> c0_n84_w173, 
            w174=> c0_n84_w174, 
            w175=> c0_n84_w175, 
            w176=> c0_n84_w176, 
            w177=> c0_n84_w177, 
            w178=> c0_n84_w178, 
            w179=> c0_n84_w179, 
            w180=> c0_n84_w180, 
            w181=> c0_n84_w181, 
            w182=> c0_n84_w182, 
            w183=> c0_n84_w183, 
            w184=> c0_n84_w184, 
            w185=> c0_n84_w185, 
            w186=> c0_n84_w186, 
            w187=> c0_n84_w187, 
            w188=> c0_n84_w188, 
            w189=> c0_n84_w189, 
            w190=> c0_n84_w190, 
            w191=> c0_n84_w191, 
            w192=> c0_n84_w192, 
            w193=> c0_n84_w193, 
            w194=> c0_n84_w194, 
            w195=> c0_n84_w195, 
            w196=> c0_n84_w196, 
            w197=> c0_n84_w197, 
            w198=> c0_n84_w198, 
            w199=> c0_n84_w199, 
            w200=> c0_n84_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n84_y
   );           
            
neuron_inst_85: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n85_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n85_w1, 
            w2=> c0_n85_w2, 
            w3=> c0_n85_w3, 
            w4=> c0_n85_w4, 
            w5=> c0_n85_w5, 
            w6=> c0_n85_w6, 
            w7=> c0_n85_w7, 
            w8=> c0_n85_w8, 
            w9=> c0_n85_w9, 
            w10=> c0_n85_w10, 
            w11=> c0_n85_w11, 
            w12=> c0_n85_w12, 
            w13=> c0_n85_w13, 
            w14=> c0_n85_w14, 
            w15=> c0_n85_w15, 
            w16=> c0_n85_w16, 
            w17=> c0_n85_w17, 
            w18=> c0_n85_w18, 
            w19=> c0_n85_w19, 
            w20=> c0_n85_w20, 
            w21=> c0_n85_w21, 
            w22=> c0_n85_w22, 
            w23=> c0_n85_w23, 
            w24=> c0_n85_w24, 
            w25=> c0_n85_w25, 
            w26=> c0_n85_w26, 
            w27=> c0_n85_w27, 
            w28=> c0_n85_w28, 
            w29=> c0_n85_w29, 
            w30=> c0_n85_w30, 
            w31=> c0_n85_w31, 
            w32=> c0_n85_w32, 
            w33=> c0_n85_w33, 
            w34=> c0_n85_w34, 
            w35=> c0_n85_w35, 
            w36=> c0_n85_w36, 
            w37=> c0_n85_w37, 
            w38=> c0_n85_w38, 
            w39=> c0_n85_w39, 
            w40=> c0_n85_w40, 
            w41=> c0_n85_w41, 
            w42=> c0_n85_w42, 
            w43=> c0_n85_w43, 
            w44=> c0_n85_w44, 
            w45=> c0_n85_w45, 
            w46=> c0_n85_w46, 
            w47=> c0_n85_w47, 
            w48=> c0_n85_w48, 
            w49=> c0_n85_w49, 
            w50=> c0_n85_w50, 
            w51=> c0_n85_w51, 
            w52=> c0_n85_w52, 
            w53=> c0_n85_w53, 
            w54=> c0_n85_w54, 
            w55=> c0_n85_w55, 
            w56=> c0_n85_w56, 
            w57=> c0_n85_w57, 
            w58=> c0_n85_w58, 
            w59=> c0_n85_w59, 
            w60=> c0_n85_w60, 
            w61=> c0_n85_w61, 
            w62=> c0_n85_w62, 
            w63=> c0_n85_w63, 
            w64=> c0_n85_w64, 
            w65=> c0_n85_w65, 
            w66=> c0_n85_w66, 
            w67=> c0_n85_w67, 
            w68=> c0_n85_w68, 
            w69=> c0_n85_w69, 
            w70=> c0_n85_w70, 
            w71=> c0_n85_w71, 
            w72=> c0_n85_w72, 
            w73=> c0_n85_w73, 
            w74=> c0_n85_w74, 
            w75=> c0_n85_w75, 
            w76=> c0_n85_w76, 
            w77=> c0_n85_w77, 
            w78=> c0_n85_w78, 
            w79=> c0_n85_w79, 
            w80=> c0_n85_w80, 
            w81=> c0_n85_w81, 
            w82=> c0_n85_w82, 
            w83=> c0_n85_w83, 
            w84=> c0_n85_w84, 
            w85=> c0_n85_w85, 
            w86=> c0_n85_w86, 
            w87=> c0_n85_w87, 
            w88=> c0_n85_w88, 
            w89=> c0_n85_w89, 
            w90=> c0_n85_w90, 
            w91=> c0_n85_w91, 
            w92=> c0_n85_w92, 
            w93=> c0_n85_w93, 
            w94=> c0_n85_w94, 
            w95=> c0_n85_w95, 
            w96=> c0_n85_w96, 
            w97=> c0_n85_w97, 
            w98=> c0_n85_w98, 
            w99=> c0_n85_w99, 
            w100=> c0_n85_w100, 
            w101=> c0_n85_w101, 
            w102=> c0_n85_w102, 
            w103=> c0_n85_w103, 
            w104=> c0_n85_w104, 
            w105=> c0_n85_w105, 
            w106=> c0_n85_w106, 
            w107=> c0_n85_w107, 
            w108=> c0_n85_w108, 
            w109=> c0_n85_w109, 
            w110=> c0_n85_w110, 
            w111=> c0_n85_w111, 
            w112=> c0_n85_w112, 
            w113=> c0_n85_w113, 
            w114=> c0_n85_w114, 
            w115=> c0_n85_w115, 
            w116=> c0_n85_w116, 
            w117=> c0_n85_w117, 
            w118=> c0_n85_w118, 
            w119=> c0_n85_w119, 
            w120=> c0_n85_w120, 
            w121=> c0_n85_w121, 
            w122=> c0_n85_w122, 
            w123=> c0_n85_w123, 
            w124=> c0_n85_w124, 
            w125=> c0_n85_w125, 
            w126=> c0_n85_w126, 
            w127=> c0_n85_w127, 
            w128=> c0_n85_w128, 
            w129=> c0_n85_w129, 
            w130=> c0_n85_w130, 
            w131=> c0_n85_w131, 
            w132=> c0_n85_w132, 
            w133=> c0_n85_w133, 
            w134=> c0_n85_w134, 
            w135=> c0_n85_w135, 
            w136=> c0_n85_w136, 
            w137=> c0_n85_w137, 
            w138=> c0_n85_w138, 
            w139=> c0_n85_w139, 
            w140=> c0_n85_w140, 
            w141=> c0_n85_w141, 
            w142=> c0_n85_w142, 
            w143=> c0_n85_w143, 
            w144=> c0_n85_w144, 
            w145=> c0_n85_w145, 
            w146=> c0_n85_w146, 
            w147=> c0_n85_w147, 
            w148=> c0_n85_w148, 
            w149=> c0_n85_w149, 
            w150=> c0_n85_w150, 
            w151=> c0_n85_w151, 
            w152=> c0_n85_w152, 
            w153=> c0_n85_w153, 
            w154=> c0_n85_w154, 
            w155=> c0_n85_w155, 
            w156=> c0_n85_w156, 
            w157=> c0_n85_w157, 
            w158=> c0_n85_w158, 
            w159=> c0_n85_w159, 
            w160=> c0_n85_w160, 
            w161=> c0_n85_w161, 
            w162=> c0_n85_w162, 
            w163=> c0_n85_w163, 
            w164=> c0_n85_w164, 
            w165=> c0_n85_w165, 
            w166=> c0_n85_w166, 
            w167=> c0_n85_w167, 
            w168=> c0_n85_w168, 
            w169=> c0_n85_w169, 
            w170=> c0_n85_w170, 
            w171=> c0_n85_w171, 
            w172=> c0_n85_w172, 
            w173=> c0_n85_w173, 
            w174=> c0_n85_w174, 
            w175=> c0_n85_w175, 
            w176=> c0_n85_w176, 
            w177=> c0_n85_w177, 
            w178=> c0_n85_w178, 
            w179=> c0_n85_w179, 
            w180=> c0_n85_w180, 
            w181=> c0_n85_w181, 
            w182=> c0_n85_w182, 
            w183=> c0_n85_w183, 
            w184=> c0_n85_w184, 
            w185=> c0_n85_w185, 
            w186=> c0_n85_w186, 
            w187=> c0_n85_w187, 
            w188=> c0_n85_w188, 
            w189=> c0_n85_w189, 
            w190=> c0_n85_w190, 
            w191=> c0_n85_w191, 
            w192=> c0_n85_w192, 
            w193=> c0_n85_w193, 
            w194=> c0_n85_w194, 
            w195=> c0_n85_w195, 
            w196=> c0_n85_w196, 
            w197=> c0_n85_w197, 
            w198=> c0_n85_w198, 
            w199=> c0_n85_w199, 
            w200=> c0_n85_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n85_y
   );           
            
neuron_inst_86: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n86_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n86_w1, 
            w2=> c0_n86_w2, 
            w3=> c0_n86_w3, 
            w4=> c0_n86_w4, 
            w5=> c0_n86_w5, 
            w6=> c0_n86_w6, 
            w7=> c0_n86_w7, 
            w8=> c0_n86_w8, 
            w9=> c0_n86_w9, 
            w10=> c0_n86_w10, 
            w11=> c0_n86_w11, 
            w12=> c0_n86_w12, 
            w13=> c0_n86_w13, 
            w14=> c0_n86_w14, 
            w15=> c0_n86_w15, 
            w16=> c0_n86_w16, 
            w17=> c0_n86_w17, 
            w18=> c0_n86_w18, 
            w19=> c0_n86_w19, 
            w20=> c0_n86_w20, 
            w21=> c0_n86_w21, 
            w22=> c0_n86_w22, 
            w23=> c0_n86_w23, 
            w24=> c0_n86_w24, 
            w25=> c0_n86_w25, 
            w26=> c0_n86_w26, 
            w27=> c0_n86_w27, 
            w28=> c0_n86_w28, 
            w29=> c0_n86_w29, 
            w30=> c0_n86_w30, 
            w31=> c0_n86_w31, 
            w32=> c0_n86_w32, 
            w33=> c0_n86_w33, 
            w34=> c0_n86_w34, 
            w35=> c0_n86_w35, 
            w36=> c0_n86_w36, 
            w37=> c0_n86_w37, 
            w38=> c0_n86_w38, 
            w39=> c0_n86_w39, 
            w40=> c0_n86_w40, 
            w41=> c0_n86_w41, 
            w42=> c0_n86_w42, 
            w43=> c0_n86_w43, 
            w44=> c0_n86_w44, 
            w45=> c0_n86_w45, 
            w46=> c0_n86_w46, 
            w47=> c0_n86_w47, 
            w48=> c0_n86_w48, 
            w49=> c0_n86_w49, 
            w50=> c0_n86_w50, 
            w51=> c0_n86_w51, 
            w52=> c0_n86_w52, 
            w53=> c0_n86_w53, 
            w54=> c0_n86_w54, 
            w55=> c0_n86_w55, 
            w56=> c0_n86_w56, 
            w57=> c0_n86_w57, 
            w58=> c0_n86_w58, 
            w59=> c0_n86_w59, 
            w60=> c0_n86_w60, 
            w61=> c0_n86_w61, 
            w62=> c0_n86_w62, 
            w63=> c0_n86_w63, 
            w64=> c0_n86_w64, 
            w65=> c0_n86_w65, 
            w66=> c0_n86_w66, 
            w67=> c0_n86_w67, 
            w68=> c0_n86_w68, 
            w69=> c0_n86_w69, 
            w70=> c0_n86_w70, 
            w71=> c0_n86_w71, 
            w72=> c0_n86_w72, 
            w73=> c0_n86_w73, 
            w74=> c0_n86_w74, 
            w75=> c0_n86_w75, 
            w76=> c0_n86_w76, 
            w77=> c0_n86_w77, 
            w78=> c0_n86_w78, 
            w79=> c0_n86_w79, 
            w80=> c0_n86_w80, 
            w81=> c0_n86_w81, 
            w82=> c0_n86_w82, 
            w83=> c0_n86_w83, 
            w84=> c0_n86_w84, 
            w85=> c0_n86_w85, 
            w86=> c0_n86_w86, 
            w87=> c0_n86_w87, 
            w88=> c0_n86_w88, 
            w89=> c0_n86_w89, 
            w90=> c0_n86_w90, 
            w91=> c0_n86_w91, 
            w92=> c0_n86_w92, 
            w93=> c0_n86_w93, 
            w94=> c0_n86_w94, 
            w95=> c0_n86_w95, 
            w96=> c0_n86_w96, 
            w97=> c0_n86_w97, 
            w98=> c0_n86_w98, 
            w99=> c0_n86_w99, 
            w100=> c0_n86_w100, 
            w101=> c0_n86_w101, 
            w102=> c0_n86_w102, 
            w103=> c0_n86_w103, 
            w104=> c0_n86_w104, 
            w105=> c0_n86_w105, 
            w106=> c0_n86_w106, 
            w107=> c0_n86_w107, 
            w108=> c0_n86_w108, 
            w109=> c0_n86_w109, 
            w110=> c0_n86_w110, 
            w111=> c0_n86_w111, 
            w112=> c0_n86_w112, 
            w113=> c0_n86_w113, 
            w114=> c0_n86_w114, 
            w115=> c0_n86_w115, 
            w116=> c0_n86_w116, 
            w117=> c0_n86_w117, 
            w118=> c0_n86_w118, 
            w119=> c0_n86_w119, 
            w120=> c0_n86_w120, 
            w121=> c0_n86_w121, 
            w122=> c0_n86_w122, 
            w123=> c0_n86_w123, 
            w124=> c0_n86_w124, 
            w125=> c0_n86_w125, 
            w126=> c0_n86_w126, 
            w127=> c0_n86_w127, 
            w128=> c0_n86_w128, 
            w129=> c0_n86_w129, 
            w130=> c0_n86_w130, 
            w131=> c0_n86_w131, 
            w132=> c0_n86_w132, 
            w133=> c0_n86_w133, 
            w134=> c0_n86_w134, 
            w135=> c0_n86_w135, 
            w136=> c0_n86_w136, 
            w137=> c0_n86_w137, 
            w138=> c0_n86_w138, 
            w139=> c0_n86_w139, 
            w140=> c0_n86_w140, 
            w141=> c0_n86_w141, 
            w142=> c0_n86_w142, 
            w143=> c0_n86_w143, 
            w144=> c0_n86_w144, 
            w145=> c0_n86_w145, 
            w146=> c0_n86_w146, 
            w147=> c0_n86_w147, 
            w148=> c0_n86_w148, 
            w149=> c0_n86_w149, 
            w150=> c0_n86_w150, 
            w151=> c0_n86_w151, 
            w152=> c0_n86_w152, 
            w153=> c0_n86_w153, 
            w154=> c0_n86_w154, 
            w155=> c0_n86_w155, 
            w156=> c0_n86_w156, 
            w157=> c0_n86_w157, 
            w158=> c0_n86_w158, 
            w159=> c0_n86_w159, 
            w160=> c0_n86_w160, 
            w161=> c0_n86_w161, 
            w162=> c0_n86_w162, 
            w163=> c0_n86_w163, 
            w164=> c0_n86_w164, 
            w165=> c0_n86_w165, 
            w166=> c0_n86_w166, 
            w167=> c0_n86_w167, 
            w168=> c0_n86_w168, 
            w169=> c0_n86_w169, 
            w170=> c0_n86_w170, 
            w171=> c0_n86_w171, 
            w172=> c0_n86_w172, 
            w173=> c0_n86_w173, 
            w174=> c0_n86_w174, 
            w175=> c0_n86_w175, 
            w176=> c0_n86_w176, 
            w177=> c0_n86_w177, 
            w178=> c0_n86_w178, 
            w179=> c0_n86_w179, 
            w180=> c0_n86_w180, 
            w181=> c0_n86_w181, 
            w182=> c0_n86_w182, 
            w183=> c0_n86_w183, 
            w184=> c0_n86_w184, 
            w185=> c0_n86_w185, 
            w186=> c0_n86_w186, 
            w187=> c0_n86_w187, 
            w188=> c0_n86_w188, 
            w189=> c0_n86_w189, 
            w190=> c0_n86_w190, 
            w191=> c0_n86_w191, 
            w192=> c0_n86_w192, 
            w193=> c0_n86_w193, 
            w194=> c0_n86_w194, 
            w195=> c0_n86_w195, 
            w196=> c0_n86_w196, 
            w197=> c0_n86_w197, 
            w198=> c0_n86_w198, 
            w199=> c0_n86_w199, 
            w200=> c0_n86_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n86_y
   );           
            
neuron_inst_87: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n87_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n87_w1, 
            w2=> c0_n87_w2, 
            w3=> c0_n87_w3, 
            w4=> c0_n87_w4, 
            w5=> c0_n87_w5, 
            w6=> c0_n87_w6, 
            w7=> c0_n87_w7, 
            w8=> c0_n87_w8, 
            w9=> c0_n87_w9, 
            w10=> c0_n87_w10, 
            w11=> c0_n87_w11, 
            w12=> c0_n87_w12, 
            w13=> c0_n87_w13, 
            w14=> c0_n87_w14, 
            w15=> c0_n87_w15, 
            w16=> c0_n87_w16, 
            w17=> c0_n87_w17, 
            w18=> c0_n87_w18, 
            w19=> c0_n87_w19, 
            w20=> c0_n87_w20, 
            w21=> c0_n87_w21, 
            w22=> c0_n87_w22, 
            w23=> c0_n87_w23, 
            w24=> c0_n87_w24, 
            w25=> c0_n87_w25, 
            w26=> c0_n87_w26, 
            w27=> c0_n87_w27, 
            w28=> c0_n87_w28, 
            w29=> c0_n87_w29, 
            w30=> c0_n87_w30, 
            w31=> c0_n87_w31, 
            w32=> c0_n87_w32, 
            w33=> c0_n87_w33, 
            w34=> c0_n87_w34, 
            w35=> c0_n87_w35, 
            w36=> c0_n87_w36, 
            w37=> c0_n87_w37, 
            w38=> c0_n87_w38, 
            w39=> c0_n87_w39, 
            w40=> c0_n87_w40, 
            w41=> c0_n87_w41, 
            w42=> c0_n87_w42, 
            w43=> c0_n87_w43, 
            w44=> c0_n87_w44, 
            w45=> c0_n87_w45, 
            w46=> c0_n87_w46, 
            w47=> c0_n87_w47, 
            w48=> c0_n87_w48, 
            w49=> c0_n87_w49, 
            w50=> c0_n87_w50, 
            w51=> c0_n87_w51, 
            w52=> c0_n87_w52, 
            w53=> c0_n87_w53, 
            w54=> c0_n87_w54, 
            w55=> c0_n87_w55, 
            w56=> c0_n87_w56, 
            w57=> c0_n87_w57, 
            w58=> c0_n87_w58, 
            w59=> c0_n87_w59, 
            w60=> c0_n87_w60, 
            w61=> c0_n87_w61, 
            w62=> c0_n87_w62, 
            w63=> c0_n87_w63, 
            w64=> c0_n87_w64, 
            w65=> c0_n87_w65, 
            w66=> c0_n87_w66, 
            w67=> c0_n87_w67, 
            w68=> c0_n87_w68, 
            w69=> c0_n87_w69, 
            w70=> c0_n87_w70, 
            w71=> c0_n87_w71, 
            w72=> c0_n87_w72, 
            w73=> c0_n87_w73, 
            w74=> c0_n87_w74, 
            w75=> c0_n87_w75, 
            w76=> c0_n87_w76, 
            w77=> c0_n87_w77, 
            w78=> c0_n87_w78, 
            w79=> c0_n87_w79, 
            w80=> c0_n87_w80, 
            w81=> c0_n87_w81, 
            w82=> c0_n87_w82, 
            w83=> c0_n87_w83, 
            w84=> c0_n87_w84, 
            w85=> c0_n87_w85, 
            w86=> c0_n87_w86, 
            w87=> c0_n87_w87, 
            w88=> c0_n87_w88, 
            w89=> c0_n87_w89, 
            w90=> c0_n87_w90, 
            w91=> c0_n87_w91, 
            w92=> c0_n87_w92, 
            w93=> c0_n87_w93, 
            w94=> c0_n87_w94, 
            w95=> c0_n87_w95, 
            w96=> c0_n87_w96, 
            w97=> c0_n87_w97, 
            w98=> c0_n87_w98, 
            w99=> c0_n87_w99, 
            w100=> c0_n87_w100, 
            w101=> c0_n87_w101, 
            w102=> c0_n87_w102, 
            w103=> c0_n87_w103, 
            w104=> c0_n87_w104, 
            w105=> c0_n87_w105, 
            w106=> c0_n87_w106, 
            w107=> c0_n87_w107, 
            w108=> c0_n87_w108, 
            w109=> c0_n87_w109, 
            w110=> c0_n87_w110, 
            w111=> c0_n87_w111, 
            w112=> c0_n87_w112, 
            w113=> c0_n87_w113, 
            w114=> c0_n87_w114, 
            w115=> c0_n87_w115, 
            w116=> c0_n87_w116, 
            w117=> c0_n87_w117, 
            w118=> c0_n87_w118, 
            w119=> c0_n87_w119, 
            w120=> c0_n87_w120, 
            w121=> c0_n87_w121, 
            w122=> c0_n87_w122, 
            w123=> c0_n87_w123, 
            w124=> c0_n87_w124, 
            w125=> c0_n87_w125, 
            w126=> c0_n87_w126, 
            w127=> c0_n87_w127, 
            w128=> c0_n87_w128, 
            w129=> c0_n87_w129, 
            w130=> c0_n87_w130, 
            w131=> c0_n87_w131, 
            w132=> c0_n87_w132, 
            w133=> c0_n87_w133, 
            w134=> c0_n87_w134, 
            w135=> c0_n87_w135, 
            w136=> c0_n87_w136, 
            w137=> c0_n87_w137, 
            w138=> c0_n87_w138, 
            w139=> c0_n87_w139, 
            w140=> c0_n87_w140, 
            w141=> c0_n87_w141, 
            w142=> c0_n87_w142, 
            w143=> c0_n87_w143, 
            w144=> c0_n87_w144, 
            w145=> c0_n87_w145, 
            w146=> c0_n87_w146, 
            w147=> c0_n87_w147, 
            w148=> c0_n87_w148, 
            w149=> c0_n87_w149, 
            w150=> c0_n87_w150, 
            w151=> c0_n87_w151, 
            w152=> c0_n87_w152, 
            w153=> c0_n87_w153, 
            w154=> c0_n87_w154, 
            w155=> c0_n87_w155, 
            w156=> c0_n87_w156, 
            w157=> c0_n87_w157, 
            w158=> c0_n87_w158, 
            w159=> c0_n87_w159, 
            w160=> c0_n87_w160, 
            w161=> c0_n87_w161, 
            w162=> c0_n87_w162, 
            w163=> c0_n87_w163, 
            w164=> c0_n87_w164, 
            w165=> c0_n87_w165, 
            w166=> c0_n87_w166, 
            w167=> c0_n87_w167, 
            w168=> c0_n87_w168, 
            w169=> c0_n87_w169, 
            w170=> c0_n87_w170, 
            w171=> c0_n87_w171, 
            w172=> c0_n87_w172, 
            w173=> c0_n87_w173, 
            w174=> c0_n87_w174, 
            w175=> c0_n87_w175, 
            w176=> c0_n87_w176, 
            w177=> c0_n87_w177, 
            w178=> c0_n87_w178, 
            w179=> c0_n87_w179, 
            w180=> c0_n87_w180, 
            w181=> c0_n87_w181, 
            w182=> c0_n87_w182, 
            w183=> c0_n87_w183, 
            w184=> c0_n87_w184, 
            w185=> c0_n87_w185, 
            w186=> c0_n87_w186, 
            w187=> c0_n87_w187, 
            w188=> c0_n87_w188, 
            w189=> c0_n87_w189, 
            w190=> c0_n87_w190, 
            w191=> c0_n87_w191, 
            w192=> c0_n87_w192, 
            w193=> c0_n87_w193, 
            w194=> c0_n87_w194, 
            w195=> c0_n87_w195, 
            w196=> c0_n87_w196, 
            w197=> c0_n87_w197, 
            w198=> c0_n87_w198, 
            w199=> c0_n87_w199, 
            w200=> c0_n87_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n87_y
   );           
            
neuron_inst_88: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n88_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n88_w1, 
            w2=> c0_n88_w2, 
            w3=> c0_n88_w3, 
            w4=> c0_n88_w4, 
            w5=> c0_n88_w5, 
            w6=> c0_n88_w6, 
            w7=> c0_n88_w7, 
            w8=> c0_n88_w8, 
            w9=> c0_n88_w9, 
            w10=> c0_n88_w10, 
            w11=> c0_n88_w11, 
            w12=> c0_n88_w12, 
            w13=> c0_n88_w13, 
            w14=> c0_n88_w14, 
            w15=> c0_n88_w15, 
            w16=> c0_n88_w16, 
            w17=> c0_n88_w17, 
            w18=> c0_n88_w18, 
            w19=> c0_n88_w19, 
            w20=> c0_n88_w20, 
            w21=> c0_n88_w21, 
            w22=> c0_n88_w22, 
            w23=> c0_n88_w23, 
            w24=> c0_n88_w24, 
            w25=> c0_n88_w25, 
            w26=> c0_n88_w26, 
            w27=> c0_n88_w27, 
            w28=> c0_n88_w28, 
            w29=> c0_n88_w29, 
            w30=> c0_n88_w30, 
            w31=> c0_n88_w31, 
            w32=> c0_n88_w32, 
            w33=> c0_n88_w33, 
            w34=> c0_n88_w34, 
            w35=> c0_n88_w35, 
            w36=> c0_n88_w36, 
            w37=> c0_n88_w37, 
            w38=> c0_n88_w38, 
            w39=> c0_n88_w39, 
            w40=> c0_n88_w40, 
            w41=> c0_n88_w41, 
            w42=> c0_n88_w42, 
            w43=> c0_n88_w43, 
            w44=> c0_n88_w44, 
            w45=> c0_n88_w45, 
            w46=> c0_n88_w46, 
            w47=> c0_n88_w47, 
            w48=> c0_n88_w48, 
            w49=> c0_n88_w49, 
            w50=> c0_n88_w50, 
            w51=> c0_n88_w51, 
            w52=> c0_n88_w52, 
            w53=> c0_n88_w53, 
            w54=> c0_n88_w54, 
            w55=> c0_n88_w55, 
            w56=> c0_n88_w56, 
            w57=> c0_n88_w57, 
            w58=> c0_n88_w58, 
            w59=> c0_n88_w59, 
            w60=> c0_n88_w60, 
            w61=> c0_n88_w61, 
            w62=> c0_n88_w62, 
            w63=> c0_n88_w63, 
            w64=> c0_n88_w64, 
            w65=> c0_n88_w65, 
            w66=> c0_n88_w66, 
            w67=> c0_n88_w67, 
            w68=> c0_n88_w68, 
            w69=> c0_n88_w69, 
            w70=> c0_n88_w70, 
            w71=> c0_n88_w71, 
            w72=> c0_n88_w72, 
            w73=> c0_n88_w73, 
            w74=> c0_n88_w74, 
            w75=> c0_n88_w75, 
            w76=> c0_n88_w76, 
            w77=> c0_n88_w77, 
            w78=> c0_n88_w78, 
            w79=> c0_n88_w79, 
            w80=> c0_n88_w80, 
            w81=> c0_n88_w81, 
            w82=> c0_n88_w82, 
            w83=> c0_n88_w83, 
            w84=> c0_n88_w84, 
            w85=> c0_n88_w85, 
            w86=> c0_n88_w86, 
            w87=> c0_n88_w87, 
            w88=> c0_n88_w88, 
            w89=> c0_n88_w89, 
            w90=> c0_n88_w90, 
            w91=> c0_n88_w91, 
            w92=> c0_n88_w92, 
            w93=> c0_n88_w93, 
            w94=> c0_n88_w94, 
            w95=> c0_n88_w95, 
            w96=> c0_n88_w96, 
            w97=> c0_n88_w97, 
            w98=> c0_n88_w98, 
            w99=> c0_n88_w99, 
            w100=> c0_n88_w100, 
            w101=> c0_n88_w101, 
            w102=> c0_n88_w102, 
            w103=> c0_n88_w103, 
            w104=> c0_n88_w104, 
            w105=> c0_n88_w105, 
            w106=> c0_n88_w106, 
            w107=> c0_n88_w107, 
            w108=> c0_n88_w108, 
            w109=> c0_n88_w109, 
            w110=> c0_n88_w110, 
            w111=> c0_n88_w111, 
            w112=> c0_n88_w112, 
            w113=> c0_n88_w113, 
            w114=> c0_n88_w114, 
            w115=> c0_n88_w115, 
            w116=> c0_n88_w116, 
            w117=> c0_n88_w117, 
            w118=> c0_n88_w118, 
            w119=> c0_n88_w119, 
            w120=> c0_n88_w120, 
            w121=> c0_n88_w121, 
            w122=> c0_n88_w122, 
            w123=> c0_n88_w123, 
            w124=> c0_n88_w124, 
            w125=> c0_n88_w125, 
            w126=> c0_n88_w126, 
            w127=> c0_n88_w127, 
            w128=> c0_n88_w128, 
            w129=> c0_n88_w129, 
            w130=> c0_n88_w130, 
            w131=> c0_n88_w131, 
            w132=> c0_n88_w132, 
            w133=> c0_n88_w133, 
            w134=> c0_n88_w134, 
            w135=> c0_n88_w135, 
            w136=> c0_n88_w136, 
            w137=> c0_n88_w137, 
            w138=> c0_n88_w138, 
            w139=> c0_n88_w139, 
            w140=> c0_n88_w140, 
            w141=> c0_n88_w141, 
            w142=> c0_n88_w142, 
            w143=> c0_n88_w143, 
            w144=> c0_n88_w144, 
            w145=> c0_n88_w145, 
            w146=> c0_n88_w146, 
            w147=> c0_n88_w147, 
            w148=> c0_n88_w148, 
            w149=> c0_n88_w149, 
            w150=> c0_n88_w150, 
            w151=> c0_n88_w151, 
            w152=> c0_n88_w152, 
            w153=> c0_n88_w153, 
            w154=> c0_n88_w154, 
            w155=> c0_n88_w155, 
            w156=> c0_n88_w156, 
            w157=> c0_n88_w157, 
            w158=> c0_n88_w158, 
            w159=> c0_n88_w159, 
            w160=> c0_n88_w160, 
            w161=> c0_n88_w161, 
            w162=> c0_n88_w162, 
            w163=> c0_n88_w163, 
            w164=> c0_n88_w164, 
            w165=> c0_n88_w165, 
            w166=> c0_n88_w166, 
            w167=> c0_n88_w167, 
            w168=> c0_n88_w168, 
            w169=> c0_n88_w169, 
            w170=> c0_n88_w170, 
            w171=> c0_n88_w171, 
            w172=> c0_n88_w172, 
            w173=> c0_n88_w173, 
            w174=> c0_n88_w174, 
            w175=> c0_n88_w175, 
            w176=> c0_n88_w176, 
            w177=> c0_n88_w177, 
            w178=> c0_n88_w178, 
            w179=> c0_n88_w179, 
            w180=> c0_n88_w180, 
            w181=> c0_n88_w181, 
            w182=> c0_n88_w182, 
            w183=> c0_n88_w183, 
            w184=> c0_n88_w184, 
            w185=> c0_n88_w185, 
            w186=> c0_n88_w186, 
            w187=> c0_n88_w187, 
            w188=> c0_n88_w188, 
            w189=> c0_n88_w189, 
            w190=> c0_n88_w190, 
            w191=> c0_n88_w191, 
            w192=> c0_n88_w192, 
            w193=> c0_n88_w193, 
            w194=> c0_n88_w194, 
            w195=> c0_n88_w195, 
            w196=> c0_n88_w196, 
            w197=> c0_n88_w197, 
            w198=> c0_n88_w198, 
            w199=> c0_n88_w199, 
            w200=> c0_n88_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n88_y
   );           
            
neuron_inst_89: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n89_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n89_w1, 
            w2=> c0_n89_w2, 
            w3=> c0_n89_w3, 
            w4=> c0_n89_w4, 
            w5=> c0_n89_w5, 
            w6=> c0_n89_w6, 
            w7=> c0_n89_w7, 
            w8=> c0_n89_w8, 
            w9=> c0_n89_w9, 
            w10=> c0_n89_w10, 
            w11=> c0_n89_w11, 
            w12=> c0_n89_w12, 
            w13=> c0_n89_w13, 
            w14=> c0_n89_w14, 
            w15=> c0_n89_w15, 
            w16=> c0_n89_w16, 
            w17=> c0_n89_w17, 
            w18=> c0_n89_w18, 
            w19=> c0_n89_w19, 
            w20=> c0_n89_w20, 
            w21=> c0_n89_w21, 
            w22=> c0_n89_w22, 
            w23=> c0_n89_w23, 
            w24=> c0_n89_w24, 
            w25=> c0_n89_w25, 
            w26=> c0_n89_w26, 
            w27=> c0_n89_w27, 
            w28=> c0_n89_w28, 
            w29=> c0_n89_w29, 
            w30=> c0_n89_w30, 
            w31=> c0_n89_w31, 
            w32=> c0_n89_w32, 
            w33=> c0_n89_w33, 
            w34=> c0_n89_w34, 
            w35=> c0_n89_w35, 
            w36=> c0_n89_w36, 
            w37=> c0_n89_w37, 
            w38=> c0_n89_w38, 
            w39=> c0_n89_w39, 
            w40=> c0_n89_w40, 
            w41=> c0_n89_w41, 
            w42=> c0_n89_w42, 
            w43=> c0_n89_w43, 
            w44=> c0_n89_w44, 
            w45=> c0_n89_w45, 
            w46=> c0_n89_w46, 
            w47=> c0_n89_w47, 
            w48=> c0_n89_w48, 
            w49=> c0_n89_w49, 
            w50=> c0_n89_w50, 
            w51=> c0_n89_w51, 
            w52=> c0_n89_w52, 
            w53=> c0_n89_w53, 
            w54=> c0_n89_w54, 
            w55=> c0_n89_w55, 
            w56=> c0_n89_w56, 
            w57=> c0_n89_w57, 
            w58=> c0_n89_w58, 
            w59=> c0_n89_w59, 
            w60=> c0_n89_w60, 
            w61=> c0_n89_w61, 
            w62=> c0_n89_w62, 
            w63=> c0_n89_w63, 
            w64=> c0_n89_w64, 
            w65=> c0_n89_w65, 
            w66=> c0_n89_w66, 
            w67=> c0_n89_w67, 
            w68=> c0_n89_w68, 
            w69=> c0_n89_w69, 
            w70=> c0_n89_w70, 
            w71=> c0_n89_w71, 
            w72=> c0_n89_w72, 
            w73=> c0_n89_w73, 
            w74=> c0_n89_w74, 
            w75=> c0_n89_w75, 
            w76=> c0_n89_w76, 
            w77=> c0_n89_w77, 
            w78=> c0_n89_w78, 
            w79=> c0_n89_w79, 
            w80=> c0_n89_w80, 
            w81=> c0_n89_w81, 
            w82=> c0_n89_w82, 
            w83=> c0_n89_w83, 
            w84=> c0_n89_w84, 
            w85=> c0_n89_w85, 
            w86=> c0_n89_w86, 
            w87=> c0_n89_w87, 
            w88=> c0_n89_w88, 
            w89=> c0_n89_w89, 
            w90=> c0_n89_w90, 
            w91=> c0_n89_w91, 
            w92=> c0_n89_w92, 
            w93=> c0_n89_w93, 
            w94=> c0_n89_w94, 
            w95=> c0_n89_w95, 
            w96=> c0_n89_w96, 
            w97=> c0_n89_w97, 
            w98=> c0_n89_w98, 
            w99=> c0_n89_w99, 
            w100=> c0_n89_w100, 
            w101=> c0_n89_w101, 
            w102=> c0_n89_w102, 
            w103=> c0_n89_w103, 
            w104=> c0_n89_w104, 
            w105=> c0_n89_w105, 
            w106=> c0_n89_w106, 
            w107=> c0_n89_w107, 
            w108=> c0_n89_w108, 
            w109=> c0_n89_w109, 
            w110=> c0_n89_w110, 
            w111=> c0_n89_w111, 
            w112=> c0_n89_w112, 
            w113=> c0_n89_w113, 
            w114=> c0_n89_w114, 
            w115=> c0_n89_w115, 
            w116=> c0_n89_w116, 
            w117=> c0_n89_w117, 
            w118=> c0_n89_w118, 
            w119=> c0_n89_w119, 
            w120=> c0_n89_w120, 
            w121=> c0_n89_w121, 
            w122=> c0_n89_w122, 
            w123=> c0_n89_w123, 
            w124=> c0_n89_w124, 
            w125=> c0_n89_w125, 
            w126=> c0_n89_w126, 
            w127=> c0_n89_w127, 
            w128=> c0_n89_w128, 
            w129=> c0_n89_w129, 
            w130=> c0_n89_w130, 
            w131=> c0_n89_w131, 
            w132=> c0_n89_w132, 
            w133=> c0_n89_w133, 
            w134=> c0_n89_w134, 
            w135=> c0_n89_w135, 
            w136=> c0_n89_w136, 
            w137=> c0_n89_w137, 
            w138=> c0_n89_w138, 
            w139=> c0_n89_w139, 
            w140=> c0_n89_w140, 
            w141=> c0_n89_w141, 
            w142=> c0_n89_w142, 
            w143=> c0_n89_w143, 
            w144=> c0_n89_w144, 
            w145=> c0_n89_w145, 
            w146=> c0_n89_w146, 
            w147=> c0_n89_w147, 
            w148=> c0_n89_w148, 
            w149=> c0_n89_w149, 
            w150=> c0_n89_w150, 
            w151=> c0_n89_w151, 
            w152=> c0_n89_w152, 
            w153=> c0_n89_w153, 
            w154=> c0_n89_w154, 
            w155=> c0_n89_w155, 
            w156=> c0_n89_w156, 
            w157=> c0_n89_w157, 
            w158=> c0_n89_w158, 
            w159=> c0_n89_w159, 
            w160=> c0_n89_w160, 
            w161=> c0_n89_w161, 
            w162=> c0_n89_w162, 
            w163=> c0_n89_w163, 
            w164=> c0_n89_w164, 
            w165=> c0_n89_w165, 
            w166=> c0_n89_w166, 
            w167=> c0_n89_w167, 
            w168=> c0_n89_w168, 
            w169=> c0_n89_w169, 
            w170=> c0_n89_w170, 
            w171=> c0_n89_w171, 
            w172=> c0_n89_w172, 
            w173=> c0_n89_w173, 
            w174=> c0_n89_w174, 
            w175=> c0_n89_w175, 
            w176=> c0_n89_w176, 
            w177=> c0_n89_w177, 
            w178=> c0_n89_w178, 
            w179=> c0_n89_w179, 
            w180=> c0_n89_w180, 
            w181=> c0_n89_w181, 
            w182=> c0_n89_w182, 
            w183=> c0_n89_w183, 
            w184=> c0_n89_w184, 
            w185=> c0_n89_w185, 
            w186=> c0_n89_w186, 
            w187=> c0_n89_w187, 
            w188=> c0_n89_w188, 
            w189=> c0_n89_w189, 
            w190=> c0_n89_w190, 
            w191=> c0_n89_w191, 
            w192=> c0_n89_w192, 
            w193=> c0_n89_w193, 
            w194=> c0_n89_w194, 
            w195=> c0_n89_w195, 
            w196=> c0_n89_w196, 
            w197=> c0_n89_w197, 
            w198=> c0_n89_w198, 
            w199=> c0_n89_w199, 
            w200=> c0_n89_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n89_y
   );           
            
neuron_inst_90: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n90_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n90_w1, 
            w2=> c0_n90_w2, 
            w3=> c0_n90_w3, 
            w4=> c0_n90_w4, 
            w5=> c0_n90_w5, 
            w6=> c0_n90_w6, 
            w7=> c0_n90_w7, 
            w8=> c0_n90_w8, 
            w9=> c0_n90_w9, 
            w10=> c0_n90_w10, 
            w11=> c0_n90_w11, 
            w12=> c0_n90_w12, 
            w13=> c0_n90_w13, 
            w14=> c0_n90_w14, 
            w15=> c0_n90_w15, 
            w16=> c0_n90_w16, 
            w17=> c0_n90_w17, 
            w18=> c0_n90_w18, 
            w19=> c0_n90_w19, 
            w20=> c0_n90_w20, 
            w21=> c0_n90_w21, 
            w22=> c0_n90_w22, 
            w23=> c0_n90_w23, 
            w24=> c0_n90_w24, 
            w25=> c0_n90_w25, 
            w26=> c0_n90_w26, 
            w27=> c0_n90_w27, 
            w28=> c0_n90_w28, 
            w29=> c0_n90_w29, 
            w30=> c0_n90_w30, 
            w31=> c0_n90_w31, 
            w32=> c0_n90_w32, 
            w33=> c0_n90_w33, 
            w34=> c0_n90_w34, 
            w35=> c0_n90_w35, 
            w36=> c0_n90_w36, 
            w37=> c0_n90_w37, 
            w38=> c0_n90_w38, 
            w39=> c0_n90_w39, 
            w40=> c0_n90_w40, 
            w41=> c0_n90_w41, 
            w42=> c0_n90_w42, 
            w43=> c0_n90_w43, 
            w44=> c0_n90_w44, 
            w45=> c0_n90_w45, 
            w46=> c0_n90_w46, 
            w47=> c0_n90_w47, 
            w48=> c0_n90_w48, 
            w49=> c0_n90_w49, 
            w50=> c0_n90_w50, 
            w51=> c0_n90_w51, 
            w52=> c0_n90_w52, 
            w53=> c0_n90_w53, 
            w54=> c0_n90_w54, 
            w55=> c0_n90_w55, 
            w56=> c0_n90_w56, 
            w57=> c0_n90_w57, 
            w58=> c0_n90_w58, 
            w59=> c0_n90_w59, 
            w60=> c0_n90_w60, 
            w61=> c0_n90_w61, 
            w62=> c0_n90_w62, 
            w63=> c0_n90_w63, 
            w64=> c0_n90_w64, 
            w65=> c0_n90_w65, 
            w66=> c0_n90_w66, 
            w67=> c0_n90_w67, 
            w68=> c0_n90_w68, 
            w69=> c0_n90_w69, 
            w70=> c0_n90_w70, 
            w71=> c0_n90_w71, 
            w72=> c0_n90_w72, 
            w73=> c0_n90_w73, 
            w74=> c0_n90_w74, 
            w75=> c0_n90_w75, 
            w76=> c0_n90_w76, 
            w77=> c0_n90_w77, 
            w78=> c0_n90_w78, 
            w79=> c0_n90_w79, 
            w80=> c0_n90_w80, 
            w81=> c0_n90_w81, 
            w82=> c0_n90_w82, 
            w83=> c0_n90_w83, 
            w84=> c0_n90_w84, 
            w85=> c0_n90_w85, 
            w86=> c0_n90_w86, 
            w87=> c0_n90_w87, 
            w88=> c0_n90_w88, 
            w89=> c0_n90_w89, 
            w90=> c0_n90_w90, 
            w91=> c0_n90_w91, 
            w92=> c0_n90_w92, 
            w93=> c0_n90_w93, 
            w94=> c0_n90_w94, 
            w95=> c0_n90_w95, 
            w96=> c0_n90_w96, 
            w97=> c0_n90_w97, 
            w98=> c0_n90_w98, 
            w99=> c0_n90_w99, 
            w100=> c0_n90_w100, 
            w101=> c0_n90_w101, 
            w102=> c0_n90_w102, 
            w103=> c0_n90_w103, 
            w104=> c0_n90_w104, 
            w105=> c0_n90_w105, 
            w106=> c0_n90_w106, 
            w107=> c0_n90_w107, 
            w108=> c0_n90_w108, 
            w109=> c0_n90_w109, 
            w110=> c0_n90_w110, 
            w111=> c0_n90_w111, 
            w112=> c0_n90_w112, 
            w113=> c0_n90_w113, 
            w114=> c0_n90_w114, 
            w115=> c0_n90_w115, 
            w116=> c0_n90_w116, 
            w117=> c0_n90_w117, 
            w118=> c0_n90_w118, 
            w119=> c0_n90_w119, 
            w120=> c0_n90_w120, 
            w121=> c0_n90_w121, 
            w122=> c0_n90_w122, 
            w123=> c0_n90_w123, 
            w124=> c0_n90_w124, 
            w125=> c0_n90_w125, 
            w126=> c0_n90_w126, 
            w127=> c0_n90_w127, 
            w128=> c0_n90_w128, 
            w129=> c0_n90_w129, 
            w130=> c0_n90_w130, 
            w131=> c0_n90_w131, 
            w132=> c0_n90_w132, 
            w133=> c0_n90_w133, 
            w134=> c0_n90_w134, 
            w135=> c0_n90_w135, 
            w136=> c0_n90_w136, 
            w137=> c0_n90_w137, 
            w138=> c0_n90_w138, 
            w139=> c0_n90_w139, 
            w140=> c0_n90_w140, 
            w141=> c0_n90_w141, 
            w142=> c0_n90_w142, 
            w143=> c0_n90_w143, 
            w144=> c0_n90_w144, 
            w145=> c0_n90_w145, 
            w146=> c0_n90_w146, 
            w147=> c0_n90_w147, 
            w148=> c0_n90_w148, 
            w149=> c0_n90_w149, 
            w150=> c0_n90_w150, 
            w151=> c0_n90_w151, 
            w152=> c0_n90_w152, 
            w153=> c0_n90_w153, 
            w154=> c0_n90_w154, 
            w155=> c0_n90_w155, 
            w156=> c0_n90_w156, 
            w157=> c0_n90_w157, 
            w158=> c0_n90_w158, 
            w159=> c0_n90_w159, 
            w160=> c0_n90_w160, 
            w161=> c0_n90_w161, 
            w162=> c0_n90_w162, 
            w163=> c0_n90_w163, 
            w164=> c0_n90_w164, 
            w165=> c0_n90_w165, 
            w166=> c0_n90_w166, 
            w167=> c0_n90_w167, 
            w168=> c0_n90_w168, 
            w169=> c0_n90_w169, 
            w170=> c0_n90_w170, 
            w171=> c0_n90_w171, 
            w172=> c0_n90_w172, 
            w173=> c0_n90_w173, 
            w174=> c0_n90_w174, 
            w175=> c0_n90_w175, 
            w176=> c0_n90_w176, 
            w177=> c0_n90_w177, 
            w178=> c0_n90_w178, 
            w179=> c0_n90_w179, 
            w180=> c0_n90_w180, 
            w181=> c0_n90_w181, 
            w182=> c0_n90_w182, 
            w183=> c0_n90_w183, 
            w184=> c0_n90_w184, 
            w185=> c0_n90_w185, 
            w186=> c0_n90_w186, 
            w187=> c0_n90_w187, 
            w188=> c0_n90_w188, 
            w189=> c0_n90_w189, 
            w190=> c0_n90_w190, 
            w191=> c0_n90_w191, 
            w192=> c0_n90_w192, 
            w193=> c0_n90_w193, 
            w194=> c0_n90_w194, 
            w195=> c0_n90_w195, 
            w196=> c0_n90_w196, 
            w197=> c0_n90_w197, 
            w198=> c0_n90_w198, 
            w199=> c0_n90_w199, 
            w200=> c0_n90_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n90_y
   );           
            
neuron_inst_91: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n91_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n91_w1, 
            w2=> c0_n91_w2, 
            w3=> c0_n91_w3, 
            w4=> c0_n91_w4, 
            w5=> c0_n91_w5, 
            w6=> c0_n91_w6, 
            w7=> c0_n91_w7, 
            w8=> c0_n91_w8, 
            w9=> c0_n91_w9, 
            w10=> c0_n91_w10, 
            w11=> c0_n91_w11, 
            w12=> c0_n91_w12, 
            w13=> c0_n91_w13, 
            w14=> c0_n91_w14, 
            w15=> c0_n91_w15, 
            w16=> c0_n91_w16, 
            w17=> c0_n91_w17, 
            w18=> c0_n91_w18, 
            w19=> c0_n91_w19, 
            w20=> c0_n91_w20, 
            w21=> c0_n91_w21, 
            w22=> c0_n91_w22, 
            w23=> c0_n91_w23, 
            w24=> c0_n91_w24, 
            w25=> c0_n91_w25, 
            w26=> c0_n91_w26, 
            w27=> c0_n91_w27, 
            w28=> c0_n91_w28, 
            w29=> c0_n91_w29, 
            w30=> c0_n91_w30, 
            w31=> c0_n91_w31, 
            w32=> c0_n91_w32, 
            w33=> c0_n91_w33, 
            w34=> c0_n91_w34, 
            w35=> c0_n91_w35, 
            w36=> c0_n91_w36, 
            w37=> c0_n91_w37, 
            w38=> c0_n91_w38, 
            w39=> c0_n91_w39, 
            w40=> c0_n91_w40, 
            w41=> c0_n91_w41, 
            w42=> c0_n91_w42, 
            w43=> c0_n91_w43, 
            w44=> c0_n91_w44, 
            w45=> c0_n91_w45, 
            w46=> c0_n91_w46, 
            w47=> c0_n91_w47, 
            w48=> c0_n91_w48, 
            w49=> c0_n91_w49, 
            w50=> c0_n91_w50, 
            w51=> c0_n91_w51, 
            w52=> c0_n91_w52, 
            w53=> c0_n91_w53, 
            w54=> c0_n91_w54, 
            w55=> c0_n91_w55, 
            w56=> c0_n91_w56, 
            w57=> c0_n91_w57, 
            w58=> c0_n91_w58, 
            w59=> c0_n91_w59, 
            w60=> c0_n91_w60, 
            w61=> c0_n91_w61, 
            w62=> c0_n91_w62, 
            w63=> c0_n91_w63, 
            w64=> c0_n91_w64, 
            w65=> c0_n91_w65, 
            w66=> c0_n91_w66, 
            w67=> c0_n91_w67, 
            w68=> c0_n91_w68, 
            w69=> c0_n91_w69, 
            w70=> c0_n91_w70, 
            w71=> c0_n91_w71, 
            w72=> c0_n91_w72, 
            w73=> c0_n91_w73, 
            w74=> c0_n91_w74, 
            w75=> c0_n91_w75, 
            w76=> c0_n91_w76, 
            w77=> c0_n91_w77, 
            w78=> c0_n91_w78, 
            w79=> c0_n91_w79, 
            w80=> c0_n91_w80, 
            w81=> c0_n91_w81, 
            w82=> c0_n91_w82, 
            w83=> c0_n91_w83, 
            w84=> c0_n91_w84, 
            w85=> c0_n91_w85, 
            w86=> c0_n91_w86, 
            w87=> c0_n91_w87, 
            w88=> c0_n91_w88, 
            w89=> c0_n91_w89, 
            w90=> c0_n91_w90, 
            w91=> c0_n91_w91, 
            w92=> c0_n91_w92, 
            w93=> c0_n91_w93, 
            w94=> c0_n91_w94, 
            w95=> c0_n91_w95, 
            w96=> c0_n91_w96, 
            w97=> c0_n91_w97, 
            w98=> c0_n91_w98, 
            w99=> c0_n91_w99, 
            w100=> c0_n91_w100, 
            w101=> c0_n91_w101, 
            w102=> c0_n91_w102, 
            w103=> c0_n91_w103, 
            w104=> c0_n91_w104, 
            w105=> c0_n91_w105, 
            w106=> c0_n91_w106, 
            w107=> c0_n91_w107, 
            w108=> c0_n91_w108, 
            w109=> c0_n91_w109, 
            w110=> c0_n91_w110, 
            w111=> c0_n91_w111, 
            w112=> c0_n91_w112, 
            w113=> c0_n91_w113, 
            w114=> c0_n91_w114, 
            w115=> c0_n91_w115, 
            w116=> c0_n91_w116, 
            w117=> c0_n91_w117, 
            w118=> c0_n91_w118, 
            w119=> c0_n91_w119, 
            w120=> c0_n91_w120, 
            w121=> c0_n91_w121, 
            w122=> c0_n91_w122, 
            w123=> c0_n91_w123, 
            w124=> c0_n91_w124, 
            w125=> c0_n91_w125, 
            w126=> c0_n91_w126, 
            w127=> c0_n91_w127, 
            w128=> c0_n91_w128, 
            w129=> c0_n91_w129, 
            w130=> c0_n91_w130, 
            w131=> c0_n91_w131, 
            w132=> c0_n91_w132, 
            w133=> c0_n91_w133, 
            w134=> c0_n91_w134, 
            w135=> c0_n91_w135, 
            w136=> c0_n91_w136, 
            w137=> c0_n91_w137, 
            w138=> c0_n91_w138, 
            w139=> c0_n91_w139, 
            w140=> c0_n91_w140, 
            w141=> c0_n91_w141, 
            w142=> c0_n91_w142, 
            w143=> c0_n91_w143, 
            w144=> c0_n91_w144, 
            w145=> c0_n91_w145, 
            w146=> c0_n91_w146, 
            w147=> c0_n91_w147, 
            w148=> c0_n91_w148, 
            w149=> c0_n91_w149, 
            w150=> c0_n91_w150, 
            w151=> c0_n91_w151, 
            w152=> c0_n91_w152, 
            w153=> c0_n91_w153, 
            w154=> c0_n91_w154, 
            w155=> c0_n91_w155, 
            w156=> c0_n91_w156, 
            w157=> c0_n91_w157, 
            w158=> c0_n91_w158, 
            w159=> c0_n91_w159, 
            w160=> c0_n91_w160, 
            w161=> c0_n91_w161, 
            w162=> c0_n91_w162, 
            w163=> c0_n91_w163, 
            w164=> c0_n91_w164, 
            w165=> c0_n91_w165, 
            w166=> c0_n91_w166, 
            w167=> c0_n91_w167, 
            w168=> c0_n91_w168, 
            w169=> c0_n91_w169, 
            w170=> c0_n91_w170, 
            w171=> c0_n91_w171, 
            w172=> c0_n91_w172, 
            w173=> c0_n91_w173, 
            w174=> c0_n91_w174, 
            w175=> c0_n91_w175, 
            w176=> c0_n91_w176, 
            w177=> c0_n91_w177, 
            w178=> c0_n91_w178, 
            w179=> c0_n91_w179, 
            w180=> c0_n91_w180, 
            w181=> c0_n91_w181, 
            w182=> c0_n91_w182, 
            w183=> c0_n91_w183, 
            w184=> c0_n91_w184, 
            w185=> c0_n91_w185, 
            w186=> c0_n91_w186, 
            w187=> c0_n91_w187, 
            w188=> c0_n91_w188, 
            w189=> c0_n91_w189, 
            w190=> c0_n91_w190, 
            w191=> c0_n91_w191, 
            w192=> c0_n91_w192, 
            w193=> c0_n91_w193, 
            w194=> c0_n91_w194, 
            w195=> c0_n91_w195, 
            w196=> c0_n91_w196, 
            w197=> c0_n91_w197, 
            w198=> c0_n91_w198, 
            w199=> c0_n91_w199, 
            w200=> c0_n91_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n91_y
   );           
            
neuron_inst_92: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n92_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n92_w1, 
            w2=> c0_n92_w2, 
            w3=> c0_n92_w3, 
            w4=> c0_n92_w4, 
            w5=> c0_n92_w5, 
            w6=> c0_n92_w6, 
            w7=> c0_n92_w7, 
            w8=> c0_n92_w8, 
            w9=> c0_n92_w9, 
            w10=> c0_n92_w10, 
            w11=> c0_n92_w11, 
            w12=> c0_n92_w12, 
            w13=> c0_n92_w13, 
            w14=> c0_n92_w14, 
            w15=> c0_n92_w15, 
            w16=> c0_n92_w16, 
            w17=> c0_n92_w17, 
            w18=> c0_n92_w18, 
            w19=> c0_n92_w19, 
            w20=> c0_n92_w20, 
            w21=> c0_n92_w21, 
            w22=> c0_n92_w22, 
            w23=> c0_n92_w23, 
            w24=> c0_n92_w24, 
            w25=> c0_n92_w25, 
            w26=> c0_n92_w26, 
            w27=> c0_n92_w27, 
            w28=> c0_n92_w28, 
            w29=> c0_n92_w29, 
            w30=> c0_n92_w30, 
            w31=> c0_n92_w31, 
            w32=> c0_n92_w32, 
            w33=> c0_n92_w33, 
            w34=> c0_n92_w34, 
            w35=> c0_n92_w35, 
            w36=> c0_n92_w36, 
            w37=> c0_n92_w37, 
            w38=> c0_n92_w38, 
            w39=> c0_n92_w39, 
            w40=> c0_n92_w40, 
            w41=> c0_n92_w41, 
            w42=> c0_n92_w42, 
            w43=> c0_n92_w43, 
            w44=> c0_n92_w44, 
            w45=> c0_n92_w45, 
            w46=> c0_n92_w46, 
            w47=> c0_n92_w47, 
            w48=> c0_n92_w48, 
            w49=> c0_n92_w49, 
            w50=> c0_n92_w50, 
            w51=> c0_n92_w51, 
            w52=> c0_n92_w52, 
            w53=> c0_n92_w53, 
            w54=> c0_n92_w54, 
            w55=> c0_n92_w55, 
            w56=> c0_n92_w56, 
            w57=> c0_n92_w57, 
            w58=> c0_n92_w58, 
            w59=> c0_n92_w59, 
            w60=> c0_n92_w60, 
            w61=> c0_n92_w61, 
            w62=> c0_n92_w62, 
            w63=> c0_n92_w63, 
            w64=> c0_n92_w64, 
            w65=> c0_n92_w65, 
            w66=> c0_n92_w66, 
            w67=> c0_n92_w67, 
            w68=> c0_n92_w68, 
            w69=> c0_n92_w69, 
            w70=> c0_n92_w70, 
            w71=> c0_n92_w71, 
            w72=> c0_n92_w72, 
            w73=> c0_n92_w73, 
            w74=> c0_n92_w74, 
            w75=> c0_n92_w75, 
            w76=> c0_n92_w76, 
            w77=> c0_n92_w77, 
            w78=> c0_n92_w78, 
            w79=> c0_n92_w79, 
            w80=> c0_n92_w80, 
            w81=> c0_n92_w81, 
            w82=> c0_n92_w82, 
            w83=> c0_n92_w83, 
            w84=> c0_n92_w84, 
            w85=> c0_n92_w85, 
            w86=> c0_n92_w86, 
            w87=> c0_n92_w87, 
            w88=> c0_n92_w88, 
            w89=> c0_n92_w89, 
            w90=> c0_n92_w90, 
            w91=> c0_n92_w91, 
            w92=> c0_n92_w92, 
            w93=> c0_n92_w93, 
            w94=> c0_n92_w94, 
            w95=> c0_n92_w95, 
            w96=> c0_n92_w96, 
            w97=> c0_n92_w97, 
            w98=> c0_n92_w98, 
            w99=> c0_n92_w99, 
            w100=> c0_n92_w100, 
            w101=> c0_n92_w101, 
            w102=> c0_n92_w102, 
            w103=> c0_n92_w103, 
            w104=> c0_n92_w104, 
            w105=> c0_n92_w105, 
            w106=> c0_n92_w106, 
            w107=> c0_n92_w107, 
            w108=> c0_n92_w108, 
            w109=> c0_n92_w109, 
            w110=> c0_n92_w110, 
            w111=> c0_n92_w111, 
            w112=> c0_n92_w112, 
            w113=> c0_n92_w113, 
            w114=> c0_n92_w114, 
            w115=> c0_n92_w115, 
            w116=> c0_n92_w116, 
            w117=> c0_n92_w117, 
            w118=> c0_n92_w118, 
            w119=> c0_n92_w119, 
            w120=> c0_n92_w120, 
            w121=> c0_n92_w121, 
            w122=> c0_n92_w122, 
            w123=> c0_n92_w123, 
            w124=> c0_n92_w124, 
            w125=> c0_n92_w125, 
            w126=> c0_n92_w126, 
            w127=> c0_n92_w127, 
            w128=> c0_n92_w128, 
            w129=> c0_n92_w129, 
            w130=> c0_n92_w130, 
            w131=> c0_n92_w131, 
            w132=> c0_n92_w132, 
            w133=> c0_n92_w133, 
            w134=> c0_n92_w134, 
            w135=> c0_n92_w135, 
            w136=> c0_n92_w136, 
            w137=> c0_n92_w137, 
            w138=> c0_n92_w138, 
            w139=> c0_n92_w139, 
            w140=> c0_n92_w140, 
            w141=> c0_n92_w141, 
            w142=> c0_n92_w142, 
            w143=> c0_n92_w143, 
            w144=> c0_n92_w144, 
            w145=> c0_n92_w145, 
            w146=> c0_n92_w146, 
            w147=> c0_n92_w147, 
            w148=> c0_n92_w148, 
            w149=> c0_n92_w149, 
            w150=> c0_n92_w150, 
            w151=> c0_n92_w151, 
            w152=> c0_n92_w152, 
            w153=> c0_n92_w153, 
            w154=> c0_n92_w154, 
            w155=> c0_n92_w155, 
            w156=> c0_n92_w156, 
            w157=> c0_n92_w157, 
            w158=> c0_n92_w158, 
            w159=> c0_n92_w159, 
            w160=> c0_n92_w160, 
            w161=> c0_n92_w161, 
            w162=> c0_n92_w162, 
            w163=> c0_n92_w163, 
            w164=> c0_n92_w164, 
            w165=> c0_n92_w165, 
            w166=> c0_n92_w166, 
            w167=> c0_n92_w167, 
            w168=> c0_n92_w168, 
            w169=> c0_n92_w169, 
            w170=> c0_n92_w170, 
            w171=> c0_n92_w171, 
            w172=> c0_n92_w172, 
            w173=> c0_n92_w173, 
            w174=> c0_n92_w174, 
            w175=> c0_n92_w175, 
            w176=> c0_n92_w176, 
            w177=> c0_n92_w177, 
            w178=> c0_n92_w178, 
            w179=> c0_n92_w179, 
            w180=> c0_n92_w180, 
            w181=> c0_n92_w181, 
            w182=> c0_n92_w182, 
            w183=> c0_n92_w183, 
            w184=> c0_n92_w184, 
            w185=> c0_n92_w185, 
            w186=> c0_n92_w186, 
            w187=> c0_n92_w187, 
            w188=> c0_n92_w188, 
            w189=> c0_n92_w189, 
            w190=> c0_n92_w190, 
            w191=> c0_n92_w191, 
            w192=> c0_n92_w192, 
            w193=> c0_n92_w193, 
            w194=> c0_n92_w194, 
            w195=> c0_n92_w195, 
            w196=> c0_n92_w196, 
            w197=> c0_n92_w197, 
            w198=> c0_n92_w198, 
            w199=> c0_n92_w199, 
            w200=> c0_n92_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n92_y
   );           
            
neuron_inst_93: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n93_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n93_w1, 
            w2=> c0_n93_w2, 
            w3=> c0_n93_w3, 
            w4=> c0_n93_w4, 
            w5=> c0_n93_w5, 
            w6=> c0_n93_w6, 
            w7=> c0_n93_w7, 
            w8=> c0_n93_w8, 
            w9=> c0_n93_w9, 
            w10=> c0_n93_w10, 
            w11=> c0_n93_w11, 
            w12=> c0_n93_w12, 
            w13=> c0_n93_w13, 
            w14=> c0_n93_w14, 
            w15=> c0_n93_w15, 
            w16=> c0_n93_w16, 
            w17=> c0_n93_w17, 
            w18=> c0_n93_w18, 
            w19=> c0_n93_w19, 
            w20=> c0_n93_w20, 
            w21=> c0_n93_w21, 
            w22=> c0_n93_w22, 
            w23=> c0_n93_w23, 
            w24=> c0_n93_w24, 
            w25=> c0_n93_w25, 
            w26=> c0_n93_w26, 
            w27=> c0_n93_w27, 
            w28=> c0_n93_w28, 
            w29=> c0_n93_w29, 
            w30=> c0_n93_w30, 
            w31=> c0_n93_w31, 
            w32=> c0_n93_w32, 
            w33=> c0_n93_w33, 
            w34=> c0_n93_w34, 
            w35=> c0_n93_w35, 
            w36=> c0_n93_w36, 
            w37=> c0_n93_w37, 
            w38=> c0_n93_w38, 
            w39=> c0_n93_w39, 
            w40=> c0_n93_w40, 
            w41=> c0_n93_w41, 
            w42=> c0_n93_w42, 
            w43=> c0_n93_w43, 
            w44=> c0_n93_w44, 
            w45=> c0_n93_w45, 
            w46=> c0_n93_w46, 
            w47=> c0_n93_w47, 
            w48=> c0_n93_w48, 
            w49=> c0_n93_w49, 
            w50=> c0_n93_w50, 
            w51=> c0_n93_w51, 
            w52=> c0_n93_w52, 
            w53=> c0_n93_w53, 
            w54=> c0_n93_w54, 
            w55=> c0_n93_w55, 
            w56=> c0_n93_w56, 
            w57=> c0_n93_w57, 
            w58=> c0_n93_w58, 
            w59=> c0_n93_w59, 
            w60=> c0_n93_w60, 
            w61=> c0_n93_w61, 
            w62=> c0_n93_w62, 
            w63=> c0_n93_w63, 
            w64=> c0_n93_w64, 
            w65=> c0_n93_w65, 
            w66=> c0_n93_w66, 
            w67=> c0_n93_w67, 
            w68=> c0_n93_w68, 
            w69=> c0_n93_w69, 
            w70=> c0_n93_w70, 
            w71=> c0_n93_w71, 
            w72=> c0_n93_w72, 
            w73=> c0_n93_w73, 
            w74=> c0_n93_w74, 
            w75=> c0_n93_w75, 
            w76=> c0_n93_w76, 
            w77=> c0_n93_w77, 
            w78=> c0_n93_w78, 
            w79=> c0_n93_w79, 
            w80=> c0_n93_w80, 
            w81=> c0_n93_w81, 
            w82=> c0_n93_w82, 
            w83=> c0_n93_w83, 
            w84=> c0_n93_w84, 
            w85=> c0_n93_w85, 
            w86=> c0_n93_w86, 
            w87=> c0_n93_w87, 
            w88=> c0_n93_w88, 
            w89=> c0_n93_w89, 
            w90=> c0_n93_w90, 
            w91=> c0_n93_w91, 
            w92=> c0_n93_w92, 
            w93=> c0_n93_w93, 
            w94=> c0_n93_w94, 
            w95=> c0_n93_w95, 
            w96=> c0_n93_w96, 
            w97=> c0_n93_w97, 
            w98=> c0_n93_w98, 
            w99=> c0_n93_w99, 
            w100=> c0_n93_w100, 
            w101=> c0_n93_w101, 
            w102=> c0_n93_w102, 
            w103=> c0_n93_w103, 
            w104=> c0_n93_w104, 
            w105=> c0_n93_w105, 
            w106=> c0_n93_w106, 
            w107=> c0_n93_w107, 
            w108=> c0_n93_w108, 
            w109=> c0_n93_w109, 
            w110=> c0_n93_w110, 
            w111=> c0_n93_w111, 
            w112=> c0_n93_w112, 
            w113=> c0_n93_w113, 
            w114=> c0_n93_w114, 
            w115=> c0_n93_w115, 
            w116=> c0_n93_w116, 
            w117=> c0_n93_w117, 
            w118=> c0_n93_w118, 
            w119=> c0_n93_w119, 
            w120=> c0_n93_w120, 
            w121=> c0_n93_w121, 
            w122=> c0_n93_w122, 
            w123=> c0_n93_w123, 
            w124=> c0_n93_w124, 
            w125=> c0_n93_w125, 
            w126=> c0_n93_w126, 
            w127=> c0_n93_w127, 
            w128=> c0_n93_w128, 
            w129=> c0_n93_w129, 
            w130=> c0_n93_w130, 
            w131=> c0_n93_w131, 
            w132=> c0_n93_w132, 
            w133=> c0_n93_w133, 
            w134=> c0_n93_w134, 
            w135=> c0_n93_w135, 
            w136=> c0_n93_w136, 
            w137=> c0_n93_w137, 
            w138=> c0_n93_w138, 
            w139=> c0_n93_w139, 
            w140=> c0_n93_w140, 
            w141=> c0_n93_w141, 
            w142=> c0_n93_w142, 
            w143=> c0_n93_w143, 
            w144=> c0_n93_w144, 
            w145=> c0_n93_w145, 
            w146=> c0_n93_w146, 
            w147=> c0_n93_w147, 
            w148=> c0_n93_w148, 
            w149=> c0_n93_w149, 
            w150=> c0_n93_w150, 
            w151=> c0_n93_w151, 
            w152=> c0_n93_w152, 
            w153=> c0_n93_w153, 
            w154=> c0_n93_w154, 
            w155=> c0_n93_w155, 
            w156=> c0_n93_w156, 
            w157=> c0_n93_w157, 
            w158=> c0_n93_w158, 
            w159=> c0_n93_w159, 
            w160=> c0_n93_w160, 
            w161=> c0_n93_w161, 
            w162=> c0_n93_w162, 
            w163=> c0_n93_w163, 
            w164=> c0_n93_w164, 
            w165=> c0_n93_w165, 
            w166=> c0_n93_w166, 
            w167=> c0_n93_w167, 
            w168=> c0_n93_w168, 
            w169=> c0_n93_w169, 
            w170=> c0_n93_w170, 
            w171=> c0_n93_w171, 
            w172=> c0_n93_w172, 
            w173=> c0_n93_w173, 
            w174=> c0_n93_w174, 
            w175=> c0_n93_w175, 
            w176=> c0_n93_w176, 
            w177=> c0_n93_w177, 
            w178=> c0_n93_w178, 
            w179=> c0_n93_w179, 
            w180=> c0_n93_w180, 
            w181=> c0_n93_w181, 
            w182=> c0_n93_w182, 
            w183=> c0_n93_w183, 
            w184=> c0_n93_w184, 
            w185=> c0_n93_w185, 
            w186=> c0_n93_w186, 
            w187=> c0_n93_w187, 
            w188=> c0_n93_w188, 
            w189=> c0_n93_w189, 
            w190=> c0_n93_w190, 
            w191=> c0_n93_w191, 
            w192=> c0_n93_w192, 
            w193=> c0_n93_w193, 
            w194=> c0_n93_w194, 
            w195=> c0_n93_w195, 
            w196=> c0_n93_w196, 
            w197=> c0_n93_w197, 
            w198=> c0_n93_w198, 
            w199=> c0_n93_w199, 
            w200=> c0_n93_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n93_y
   );           
            
neuron_inst_94: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n94_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n94_w1, 
            w2=> c0_n94_w2, 
            w3=> c0_n94_w3, 
            w4=> c0_n94_w4, 
            w5=> c0_n94_w5, 
            w6=> c0_n94_w6, 
            w7=> c0_n94_w7, 
            w8=> c0_n94_w8, 
            w9=> c0_n94_w9, 
            w10=> c0_n94_w10, 
            w11=> c0_n94_w11, 
            w12=> c0_n94_w12, 
            w13=> c0_n94_w13, 
            w14=> c0_n94_w14, 
            w15=> c0_n94_w15, 
            w16=> c0_n94_w16, 
            w17=> c0_n94_w17, 
            w18=> c0_n94_w18, 
            w19=> c0_n94_w19, 
            w20=> c0_n94_w20, 
            w21=> c0_n94_w21, 
            w22=> c0_n94_w22, 
            w23=> c0_n94_w23, 
            w24=> c0_n94_w24, 
            w25=> c0_n94_w25, 
            w26=> c0_n94_w26, 
            w27=> c0_n94_w27, 
            w28=> c0_n94_w28, 
            w29=> c0_n94_w29, 
            w30=> c0_n94_w30, 
            w31=> c0_n94_w31, 
            w32=> c0_n94_w32, 
            w33=> c0_n94_w33, 
            w34=> c0_n94_w34, 
            w35=> c0_n94_w35, 
            w36=> c0_n94_w36, 
            w37=> c0_n94_w37, 
            w38=> c0_n94_w38, 
            w39=> c0_n94_w39, 
            w40=> c0_n94_w40, 
            w41=> c0_n94_w41, 
            w42=> c0_n94_w42, 
            w43=> c0_n94_w43, 
            w44=> c0_n94_w44, 
            w45=> c0_n94_w45, 
            w46=> c0_n94_w46, 
            w47=> c0_n94_w47, 
            w48=> c0_n94_w48, 
            w49=> c0_n94_w49, 
            w50=> c0_n94_w50, 
            w51=> c0_n94_w51, 
            w52=> c0_n94_w52, 
            w53=> c0_n94_w53, 
            w54=> c0_n94_w54, 
            w55=> c0_n94_w55, 
            w56=> c0_n94_w56, 
            w57=> c0_n94_w57, 
            w58=> c0_n94_w58, 
            w59=> c0_n94_w59, 
            w60=> c0_n94_w60, 
            w61=> c0_n94_w61, 
            w62=> c0_n94_w62, 
            w63=> c0_n94_w63, 
            w64=> c0_n94_w64, 
            w65=> c0_n94_w65, 
            w66=> c0_n94_w66, 
            w67=> c0_n94_w67, 
            w68=> c0_n94_w68, 
            w69=> c0_n94_w69, 
            w70=> c0_n94_w70, 
            w71=> c0_n94_w71, 
            w72=> c0_n94_w72, 
            w73=> c0_n94_w73, 
            w74=> c0_n94_w74, 
            w75=> c0_n94_w75, 
            w76=> c0_n94_w76, 
            w77=> c0_n94_w77, 
            w78=> c0_n94_w78, 
            w79=> c0_n94_w79, 
            w80=> c0_n94_w80, 
            w81=> c0_n94_w81, 
            w82=> c0_n94_w82, 
            w83=> c0_n94_w83, 
            w84=> c0_n94_w84, 
            w85=> c0_n94_w85, 
            w86=> c0_n94_w86, 
            w87=> c0_n94_w87, 
            w88=> c0_n94_w88, 
            w89=> c0_n94_w89, 
            w90=> c0_n94_w90, 
            w91=> c0_n94_w91, 
            w92=> c0_n94_w92, 
            w93=> c0_n94_w93, 
            w94=> c0_n94_w94, 
            w95=> c0_n94_w95, 
            w96=> c0_n94_w96, 
            w97=> c0_n94_w97, 
            w98=> c0_n94_w98, 
            w99=> c0_n94_w99, 
            w100=> c0_n94_w100, 
            w101=> c0_n94_w101, 
            w102=> c0_n94_w102, 
            w103=> c0_n94_w103, 
            w104=> c0_n94_w104, 
            w105=> c0_n94_w105, 
            w106=> c0_n94_w106, 
            w107=> c0_n94_w107, 
            w108=> c0_n94_w108, 
            w109=> c0_n94_w109, 
            w110=> c0_n94_w110, 
            w111=> c0_n94_w111, 
            w112=> c0_n94_w112, 
            w113=> c0_n94_w113, 
            w114=> c0_n94_w114, 
            w115=> c0_n94_w115, 
            w116=> c0_n94_w116, 
            w117=> c0_n94_w117, 
            w118=> c0_n94_w118, 
            w119=> c0_n94_w119, 
            w120=> c0_n94_w120, 
            w121=> c0_n94_w121, 
            w122=> c0_n94_w122, 
            w123=> c0_n94_w123, 
            w124=> c0_n94_w124, 
            w125=> c0_n94_w125, 
            w126=> c0_n94_w126, 
            w127=> c0_n94_w127, 
            w128=> c0_n94_w128, 
            w129=> c0_n94_w129, 
            w130=> c0_n94_w130, 
            w131=> c0_n94_w131, 
            w132=> c0_n94_w132, 
            w133=> c0_n94_w133, 
            w134=> c0_n94_w134, 
            w135=> c0_n94_w135, 
            w136=> c0_n94_w136, 
            w137=> c0_n94_w137, 
            w138=> c0_n94_w138, 
            w139=> c0_n94_w139, 
            w140=> c0_n94_w140, 
            w141=> c0_n94_w141, 
            w142=> c0_n94_w142, 
            w143=> c0_n94_w143, 
            w144=> c0_n94_w144, 
            w145=> c0_n94_w145, 
            w146=> c0_n94_w146, 
            w147=> c0_n94_w147, 
            w148=> c0_n94_w148, 
            w149=> c0_n94_w149, 
            w150=> c0_n94_w150, 
            w151=> c0_n94_w151, 
            w152=> c0_n94_w152, 
            w153=> c0_n94_w153, 
            w154=> c0_n94_w154, 
            w155=> c0_n94_w155, 
            w156=> c0_n94_w156, 
            w157=> c0_n94_w157, 
            w158=> c0_n94_w158, 
            w159=> c0_n94_w159, 
            w160=> c0_n94_w160, 
            w161=> c0_n94_w161, 
            w162=> c0_n94_w162, 
            w163=> c0_n94_w163, 
            w164=> c0_n94_w164, 
            w165=> c0_n94_w165, 
            w166=> c0_n94_w166, 
            w167=> c0_n94_w167, 
            w168=> c0_n94_w168, 
            w169=> c0_n94_w169, 
            w170=> c0_n94_w170, 
            w171=> c0_n94_w171, 
            w172=> c0_n94_w172, 
            w173=> c0_n94_w173, 
            w174=> c0_n94_w174, 
            w175=> c0_n94_w175, 
            w176=> c0_n94_w176, 
            w177=> c0_n94_w177, 
            w178=> c0_n94_w178, 
            w179=> c0_n94_w179, 
            w180=> c0_n94_w180, 
            w181=> c0_n94_w181, 
            w182=> c0_n94_w182, 
            w183=> c0_n94_w183, 
            w184=> c0_n94_w184, 
            w185=> c0_n94_w185, 
            w186=> c0_n94_w186, 
            w187=> c0_n94_w187, 
            w188=> c0_n94_w188, 
            w189=> c0_n94_w189, 
            w190=> c0_n94_w190, 
            w191=> c0_n94_w191, 
            w192=> c0_n94_w192, 
            w193=> c0_n94_w193, 
            w194=> c0_n94_w194, 
            w195=> c0_n94_w195, 
            w196=> c0_n94_w196, 
            w197=> c0_n94_w197, 
            w198=> c0_n94_w198, 
            w199=> c0_n94_w199, 
            w200=> c0_n94_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n94_y
   );           
            
neuron_inst_95: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n95_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n95_w1, 
            w2=> c0_n95_w2, 
            w3=> c0_n95_w3, 
            w4=> c0_n95_w4, 
            w5=> c0_n95_w5, 
            w6=> c0_n95_w6, 
            w7=> c0_n95_w7, 
            w8=> c0_n95_w8, 
            w9=> c0_n95_w9, 
            w10=> c0_n95_w10, 
            w11=> c0_n95_w11, 
            w12=> c0_n95_w12, 
            w13=> c0_n95_w13, 
            w14=> c0_n95_w14, 
            w15=> c0_n95_w15, 
            w16=> c0_n95_w16, 
            w17=> c0_n95_w17, 
            w18=> c0_n95_w18, 
            w19=> c0_n95_w19, 
            w20=> c0_n95_w20, 
            w21=> c0_n95_w21, 
            w22=> c0_n95_w22, 
            w23=> c0_n95_w23, 
            w24=> c0_n95_w24, 
            w25=> c0_n95_w25, 
            w26=> c0_n95_w26, 
            w27=> c0_n95_w27, 
            w28=> c0_n95_w28, 
            w29=> c0_n95_w29, 
            w30=> c0_n95_w30, 
            w31=> c0_n95_w31, 
            w32=> c0_n95_w32, 
            w33=> c0_n95_w33, 
            w34=> c0_n95_w34, 
            w35=> c0_n95_w35, 
            w36=> c0_n95_w36, 
            w37=> c0_n95_w37, 
            w38=> c0_n95_w38, 
            w39=> c0_n95_w39, 
            w40=> c0_n95_w40, 
            w41=> c0_n95_w41, 
            w42=> c0_n95_w42, 
            w43=> c0_n95_w43, 
            w44=> c0_n95_w44, 
            w45=> c0_n95_w45, 
            w46=> c0_n95_w46, 
            w47=> c0_n95_w47, 
            w48=> c0_n95_w48, 
            w49=> c0_n95_w49, 
            w50=> c0_n95_w50, 
            w51=> c0_n95_w51, 
            w52=> c0_n95_w52, 
            w53=> c0_n95_w53, 
            w54=> c0_n95_w54, 
            w55=> c0_n95_w55, 
            w56=> c0_n95_w56, 
            w57=> c0_n95_w57, 
            w58=> c0_n95_w58, 
            w59=> c0_n95_w59, 
            w60=> c0_n95_w60, 
            w61=> c0_n95_w61, 
            w62=> c0_n95_w62, 
            w63=> c0_n95_w63, 
            w64=> c0_n95_w64, 
            w65=> c0_n95_w65, 
            w66=> c0_n95_w66, 
            w67=> c0_n95_w67, 
            w68=> c0_n95_w68, 
            w69=> c0_n95_w69, 
            w70=> c0_n95_w70, 
            w71=> c0_n95_w71, 
            w72=> c0_n95_w72, 
            w73=> c0_n95_w73, 
            w74=> c0_n95_w74, 
            w75=> c0_n95_w75, 
            w76=> c0_n95_w76, 
            w77=> c0_n95_w77, 
            w78=> c0_n95_w78, 
            w79=> c0_n95_w79, 
            w80=> c0_n95_w80, 
            w81=> c0_n95_w81, 
            w82=> c0_n95_w82, 
            w83=> c0_n95_w83, 
            w84=> c0_n95_w84, 
            w85=> c0_n95_w85, 
            w86=> c0_n95_w86, 
            w87=> c0_n95_w87, 
            w88=> c0_n95_w88, 
            w89=> c0_n95_w89, 
            w90=> c0_n95_w90, 
            w91=> c0_n95_w91, 
            w92=> c0_n95_w92, 
            w93=> c0_n95_w93, 
            w94=> c0_n95_w94, 
            w95=> c0_n95_w95, 
            w96=> c0_n95_w96, 
            w97=> c0_n95_w97, 
            w98=> c0_n95_w98, 
            w99=> c0_n95_w99, 
            w100=> c0_n95_w100, 
            w101=> c0_n95_w101, 
            w102=> c0_n95_w102, 
            w103=> c0_n95_w103, 
            w104=> c0_n95_w104, 
            w105=> c0_n95_w105, 
            w106=> c0_n95_w106, 
            w107=> c0_n95_w107, 
            w108=> c0_n95_w108, 
            w109=> c0_n95_w109, 
            w110=> c0_n95_w110, 
            w111=> c0_n95_w111, 
            w112=> c0_n95_w112, 
            w113=> c0_n95_w113, 
            w114=> c0_n95_w114, 
            w115=> c0_n95_w115, 
            w116=> c0_n95_w116, 
            w117=> c0_n95_w117, 
            w118=> c0_n95_w118, 
            w119=> c0_n95_w119, 
            w120=> c0_n95_w120, 
            w121=> c0_n95_w121, 
            w122=> c0_n95_w122, 
            w123=> c0_n95_w123, 
            w124=> c0_n95_w124, 
            w125=> c0_n95_w125, 
            w126=> c0_n95_w126, 
            w127=> c0_n95_w127, 
            w128=> c0_n95_w128, 
            w129=> c0_n95_w129, 
            w130=> c0_n95_w130, 
            w131=> c0_n95_w131, 
            w132=> c0_n95_w132, 
            w133=> c0_n95_w133, 
            w134=> c0_n95_w134, 
            w135=> c0_n95_w135, 
            w136=> c0_n95_w136, 
            w137=> c0_n95_w137, 
            w138=> c0_n95_w138, 
            w139=> c0_n95_w139, 
            w140=> c0_n95_w140, 
            w141=> c0_n95_w141, 
            w142=> c0_n95_w142, 
            w143=> c0_n95_w143, 
            w144=> c0_n95_w144, 
            w145=> c0_n95_w145, 
            w146=> c0_n95_w146, 
            w147=> c0_n95_w147, 
            w148=> c0_n95_w148, 
            w149=> c0_n95_w149, 
            w150=> c0_n95_w150, 
            w151=> c0_n95_w151, 
            w152=> c0_n95_w152, 
            w153=> c0_n95_w153, 
            w154=> c0_n95_w154, 
            w155=> c0_n95_w155, 
            w156=> c0_n95_w156, 
            w157=> c0_n95_w157, 
            w158=> c0_n95_w158, 
            w159=> c0_n95_w159, 
            w160=> c0_n95_w160, 
            w161=> c0_n95_w161, 
            w162=> c0_n95_w162, 
            w163=> c0_n95_w163, 
            w164=> c0_n95_w164, 
            w165=> c0_n95_w165, 
            w166=> c0_n95_w166, 
            w167=> c0_n95_w167, 
            w168=> c0_n95_w168, 
            w169=> c0_n95_w169, 
            w170=> c0_n95_w170, 
            w171=> c0_n95_w171, 
            w172=> c0_n95_w172, 
            w173=> c0_n95_w173, 
            w174=> c0_n95_w174, 
            w175=> c0_n95_w175, 
            w176=> c0_n95_w176, 
            w177=> c0_n95_w177, 
            w178=> c0_n95_w178, 
            w179=> c0_n95_w179, 
            w180=> c0_n95_w180, 
            w181=> c0_n95_w181, 
            w182=> c0_n95_w182, 
            w183=> c0_n95_w183, 
            w184=> c0_n95_w184, 
            w185=> c0_n95_w185, 
            w186=> c0_n95_w186, 
            w187=> c0_n95_w187, 
            w188=> c0_n95_w188, 
            w189=> c0_n95_w189, 
            w190=> c0_n95_w190, 
            w191=> c0_n95_w191, 
            w192=> c0_n95_w192, 
            w193=> c0_n95_w193, 
            w194=> c0_n95_w194, 
            w195=> c0_n95_w195, 
            w196=> c0_n95_w196, 
            w197=> c0_n95_w197, 
            w198=> c0_n95_w198, 
            w199=> c0_n95_w199, 
            w200=> c0_n95_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n95_y
   );           
            
neuron_inst_96: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n96_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n96_w1, 
            w2=> c0_n96_w2, 
            w3=> c0_n96_w3, 
            w4=> c0_n96_w4, 
            w5=> c0_n96_w5, 
            w6=> c0_n96_w6, 
            w7=> c0_n96_w7, 
            w8=> c0_n96_w8, 
            w9=> c0_n96_w9, 
            w10=> c0_n96_w10, 
            w11=> c0_n96_w11, 
            w12=> c0_n96_w12, 
            w13=> c0_n96_w13, 
            w14=> c0_n96_w14, 
            w15=> c0_n96_w15, 
            w16=> c0_n96_w16, 
            w17=> c0_n96_w17, 
            w18=> c0_n96_w18, 
            w19=> c0_n96_w19, 
            w20=> c0_n96_w20, 
            w21=> c0_n96_w21, 
            w22=> c0_n96_w22, 
            w23=> c0_n96_w23, 
            w24=> c0_n96_w24, 
            w25=> c0_n96_w25, 
            w26=> c0_n96_w26, 
            w27=> c0_n96_w27, 
            w28=> c0_n96_w28, 
            w29=> c0_n96_w29, 
            w30=> c0_n96_w30, 
            w31=> c0_n96_w31, 
            w32=> c0_n96_w32, 
            w33=> c0_n96_w33, 
            w34=> c0_n96_w34, 
            w35=> c0_n96_w35, 
            w36=> c0_n96_w36, 
            w37=> c0_n96_w37, 
            w38=> c0_n96_w38, 
            w39=> c0_n96_w39, 
            w40=> c0_n96_w40, 
            w41=> c0_n96_w41, 
            w42=> c0_n96_w42, 
            w43=> c0_n96_w43, 
            w44=> c0_n96_w44, 
            w45=> c0_n96_w45, 
            w46=> c0_n96_w46, 
            w47=> c0_n96_w47, 
            w48=> c0_n96_w48, 
            w49=> c0_n96_w49, 
            w50=> c0_n96_w50, 
            w51=> c0_n96_w51, 
            w52=> c0_n96_w52, 
            w53=> c0_n96_w53, 
            w54=> c0_n96_w54, 
            w55=> c0_n96_w55, 
            w56=> c0_n96_w56, 
            w57=> c0_n96_w57, 
            w58=> c0_n96_w58, 
            w59=> c0_n96_w59, 
            w60=> c0_n96_w60, 
            w61=> c0_n96_w61, 
            w62=> c0_n96_w62, 
            w63=> c0_n96_w63, 
            w64=> c0_n96_w64, 
            w65=> c0_n96_w65, 
            w66=> c0_n96_w66, 
            w67=> c0_n96_w67, 
            w68=> c0_n96_w68, 
            w69=> c0_n96_w69, 
            w70=> c0_n96_w70, 
            w71=> c0_n96_w71, 
            w72=> c0_n96_w72, 
            w73=> c0_n96_w73, 
            w74=> c0_n96_w74, 
            w75=> c0_n96_w75, 
            w76=> c0_n96_w76, 
            w77=> c0_n96_w77, 
            w78=> c0_n96_w78, 
            w79=> c0_n96_w79, 
            w80=> c0_n96_w80, 
            w81=> c0_n96_w81, 
            w82=> c0_n96_w82, 
            w83=> c0_n96_w83, 
            w84=> c0_n96_w84, 
            w85=> c0_n96_w85, 
            w86=> c0_n96_w86, 
            w87=> c0_n96_w87, 
            w88=> c0_n96_w88, 
            w89=> c0_n96_w89, 
            w90=> c0_n96_w90, 
            w91=> c0_n96_w91, 
            w92=> c0_n96_w92, 
            w93=> c0_n96_w93, 
            w94=> c0_n96_w94, 
            w95=> c0_n96_w95, 
            w96=> c0_n96_w96, 
            w97=> c0_n96_w97, 
            w98=> c0_n96_w98, 
            w99=> c0_n96_w99, 
            w100=> c0_n96_w100, 
            w101=> c0_n96_w101, 
            w102=> c0_n96_w102, 
            w103=> c0_n96_w103, 
            w104=> c0_n96_w104, 
            w105=> c0_n96_w105, 
            w106=> c0_n96_w106, 
            w107=> c0_n96_w107, 
            w108=> c0_n96_w108, 
            w109=> c0_n96_w109, 
            w110=> c0_n96_w110, 
            w111=> c0_n96_w111, 
            w112=> c0_n96_w112, 
            w113=> c0_n96_w113, 
            w114=> c0_n96_w114, 
            w115=> c0_n96_w115, 
            w116=> c0_n96_w116, 
            w117=> c0_n96_w117, 
            w118=> c0_n96_w118, 
            w119=> c0_n96_w119, 
            w120=> c0_n96_w120, 
            w121=> c0_n96_w121, 
            w122=> c0_n96_w122, 
            w123=> c0_n96_w123, 
            w124=> c0_n96_w124, 
            w125=> c0_n96_w125, 
            w126=> c0_n96_w126, 
            w127=> c0_n96_w127, 
            w128=> c0_n96_w128, 
            w129=> c0_n96_w129, 
            w130=> c0_n96_w130, 
            w131=> c0_n96_w131, 
            w132=> c0_n96_w132, 
            w133=> c0_n96_w133, 
            w134=> c0_n96_w134, 
            w135=> c0_n96_w135, 
            w136=> c0_n96_w136, 
            w137=> c0_n96_w137, 
            w138=> c0_n96_w138, 
            w139=> c0_n96_w139, 
            w140=> c0_n96_w140, 
            w141=> c0_n96_w141, 
            w142=> c0_n96_w142, 
            w143=> c0_n96_w143, 
            w144=> c0_n96_w144, 
            w145=> c0_n96_w145, 
            w146=> c0_n96_w146, 
            w147=> c0_n96_w147, 
            w148=> c0_n96_w148, 
            w149=> c0_n96_w149, 
            w150=> c0_n96_w150, 
            w151=> c0_n96_w151, 
            w152=> c0_n96_w152, 
            w153=> c0_n96_w153, 
            w154=> c0_n96_w154, 
            w155=> c0_n96_w155, 
            w156=> c0_n96_w156, 
            w157=> c0_n96_w157, 
            w158=> c0_n96_w158, 
            w159=> c0_n96_w159, 
            w160=> c0_n96_w160, 
            w161=> c0_n96_w161, 
            w162=> c0_n96_w162, 
            w163=> c0_n96_w163, 
            w164=> c0_n96_w164, 
            w165=> c0_n96_w165, 
            w166=> c0_n96_w166, 
            w167=> c0_n96_w167, 
            w168=> c0_n96_w168, 
            w169=> c0_n96_w169, 
            w170=> c0_n96_w170, 
            w171=> c0_n96_w171, 
            w172=> c0_n96_w172, 
            w173=> c0_n96_w173, 
            w174=> c0_n96_w174, 
            w175=> c0_n96_w175, 
            w176=> c0_n96_w176, 
            w177=> c0_n96_w177, 
            w178=> c0_n96_w178, 
            w179=> c0_n96_w179, 
            w180=> c0_n96_w180, 
            w181=> c0_n96_w181, 
            w182=> c0_n96_w182, 
            w183=> c0_n96_w183, 
            w184=> c0_n96_w184, 
            w185=> c0_n96_w185, 
            w186=> c0_n96_w186, 
            w187=> c0_n96_w187, 
            w188=> c0_n96_w188, 
            w189=> c0_n96_w189, 
            w190=> c0_n96_w190, 
            w191=> c0_n96_w191, 
            w192=> c0_n96_w192, 
            w193=> c0_n96_w193, 
            w194=> c0_n96_w194, 
            w195=> c0_n96_w195, 
            w196=> c0_n96_w196, 
            w197=> c0_n96_w197, 
            w198=> c0_n96_w198, 
            w199=> c0_n96_w199, 
            w200=> c0_n96_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n96_y
   );           
            
neuron_inst_97: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n97_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n97_w1, 
            w2=> c0_n97_w2, 
            w3=> c0_n97_w3, 
            w4=> c0_n97_w4, 
            w5=> c0_n97_w5, 
            w6=> c0_n97_w6, 
            w7=> c0_n97_w7, 
            w8=> c0_n97_w8, 
            w9=> c0_n97_w9, 
            w10=> c0_n97_w10, 
            w11=> c0_n97_w11, 
            w12=> c0_n97_w12, 
            w13=> c0_n97_w13, 
            w14=> c0_n97_w14, 
            w15=> c0_n97_w15, 
            w16=> c0_n97_w16, 
            w17=> c0_n97_w17, 
            w18=> c0_n97_w18, 
            w19=> c0_n97_w19, 
            w20=> c0_n97_w20, 
            w21=> c0_n97_w21, 
            w22=> c0_n97_w22, 
            w23=> c0_n97_w23, 
            w24=> c0_n97_w24, 
            w25=> c0_n97_w25, 
            w26=> c0_n97_w26, 
            w27=> c0_n97_w27, 
            w28=> c0_n97_w28, 
            w29=> c0_n97_w29, 
            w30=> c0_n97_w30, 
            w31=> c0_n97_w31, 
            w32=> c0_n97_w32, 
            w33=> c0_n97_w33, 
            w34=> c0_n97_w34, 
            w35=> c0_n97_w35, 
            w36=> c0_n97_w36, 
            w37=> c0_n97_w37, 
            w38=> c0_n97_w38, 
            w39=> c0_n97_w39, 
            w40=> c0_n97_w40, 
            w41=> c0_n97_w41, 
            w42=> c0_n97_w42, 
            w43=> c0_n97_w43, 
            w44=> c0_n97_w44, 
            w45=> c0_n97_w45, 
            w46=> c0_n97_w46, 
            w47=> c0_n97_w47, 
            w48=> c0_n97_w48, 
            w49=> c0_n97_w49, 
            w50=> c0_n97_w50, 
            w51=> c0_n97_w51, 
            w52=> c0_n97_w52, 
            w53=> c0_n97_w53, 
            w54=> c0_n97_w54, 
            w55=> c0_n97_w55, 
            w56=> c0_n97_w56, 
            w57=> c0_n97_w57, 
            w58=> c0_n97_w58, 
            w59=> c0_n97_w59, 
            w60=> c0_n97_w60, 
            w61=> c0_n97_w61, 
            w62=> c0_n97_w62, 
            w63=> c0_n97_w63, 
            w64=> c0_n97_w64, 
            w65=> c0_n97_w65, 
            w66=> c0_n97_w66, 
            w67=> c0_n97_w67, 
            w68=> c0_n97_w68, 
            w69=> c0_n97_w69, 
            w70=> c0_n97_w70, 
            w71=> c0_n97_w71, 
            w72=> c0_n97_w72, 
            w73=> c0_n97_w73, 
            w74=> c0_n97_w74, 
            w75=> c0_n97_w75, 
            w76=> c0_n97_w76, 
            w77=> c0_n97_w77, 
            w78=> c0_n97_w78, 
            w79=> c0_n97_w79, 
            w80=> c0_n97_w80, 
            w81=> c0_n97_w81, 
            w82=> c0_n97_w82, 
            w83=> c0_n97_w83, 
            w84=> c0_n97_w84, 
            w85=> c0_n97_w85, 
            w86=> c0_n97_w86, 
            w87=> c0_n97_w87, 
            w88=> c0_n97_w88, 
            w89=> c0_n97_w89, 
            w90=> c0_n97_w90, 
            w91=> c0_n97_w91, 
            w92=> c0_n97_w92, 
            w93=> c0_n97_w93, 
            w94=> c0_n97_w94, 
            w95=> c0_n97_w95, 
            w96=> c0_n97_w96, 
            w97=> c0_n97_w97, 
            w98=> c0_n97_w98, 
            w99=> c0_n97_w99, 
            w100=> c0_n97_w100, 
            w101=> c0_n97_w101, 
            w102=> c0_n97_w102, 
            w103=> c0_n97_w103, 
            w104=> c0_n97_w104, 
            w105=> c0_n97_w105, 
            w106=> c0_n97_w106, 
            w107=> c0_n97_w107, 
            w108=> c0_n97_w108, 
            w109=> c0_n97_w109, 
            w110=> c0_n97_w110, 
            w111=> c0_n97_w111, 
            w112=> c0_n97_w112, 
            w113=> c0_n97_w113, 
            w114=> c0_n97_w114, 
            w115=> c0_n97_w115, 
            w116=> c0_n97_w116, 
            w117=> c0_n97_w117, 
            w118=> c0_n97_w118, 
            w119=> c0_n97_w119, 
            w120=> c0_n97_w120, 
            w121=> c0_n97_w121, 
            w122=> c0_n97_w122, 
            w123=> c0_n97_w123, 
            w124=> c0_n97_w124, 
            w125=> c0_n97_w125, 
            w126=> c0_n97_w126, 
            w127=> c0_n97_w127, 
            w128=> c0_n97_w128, 
            w129=> c0_n97_w129, 
            w130=> c0_n97_w130, 
            w131=> c0_n97_w131, 
            w132=> c0_n97_w132, 
            w133=> c0_n97_w133, 
            w134=> c0_n97_w134, 
            w135=> c0_n97_w135, 
            w136=> c0_n97_w136, 
            w137=> c0_n97_w137, 
            w138=> c0_n97_w138, 
            w139=> c0_n97_w139, 
            w140=> c0_n97_w140, 
            w141=> c0_n97_w141, 
            w142=> c0_n97_w142, 
            w143=> c0_n97_w143, 
            w144=> c0_n97_w144, 
            w145=> c0_n97_w145, 
            w146=> c0_n97_w146, 
            w147=> c0_n97_w147, 
            w148=> c0_n97_w148, 
            w149=> c0_n97_w149, 
            w150=> c0_n97_w150, 
            w151=> c0_n97_w151, 
            w152=> c0_n97_w152, 
            w153=> c0_n97_w153, 
            w154=> c0_n97_w154, 
            w155=> c0_n97_w155, 
            w156=> c0_n97_w156, 
            w157=> c0_n97_w157, 
            w158=> c0_n97_w158, 
            w159=> c0_n97_w159, 
            w160=> c0_n97_w160, 
            w161=> c0_n97_w161, 
            w162=> c0_n97_w162, 
            w163=> c0_n97_w163, 
            w164=> c0_n97_w164, 
            w165=> c0_n97_w165, 
            w166=> c0_n97_w166, 
            w167=> c0_n97_w167, 
            w168=> c0_n97_w168, 
            w169=> c0_n97_w169, 
            w170=> c0_n97_w170, 
            w171=> c0_n97_w171, 
            w172=> c0_n97_w172, 
            w173=> c0_n97_w173, 
            w174=> c0_n97_w174, 
            w175=> c0_n97_w175, 
            w176=> c0_n97_w176, 
            w177=> c0_n97_w177, 
            w178=> c0_n97_w178, 
            w179=> c0_n97_w179, 
            w180=> c0_n97_w180, 
            w181=> c0_n97_w181, 
            w182=> c0_n97_w182, 
            w183=> c0_n97_w183, 
            w184=> c0_n97_w184, 
            w185=> c0_n97_w185, 
            w186=> c0_n97_w186, 
            w187=> c0_n97_w187, 
            w188=> c0_n97_w188, 
            w189=> c0_n97_w189, 
            w190=> c0_n97_w190, 
            w191=> c0_n97_w191, 
            w192=> c0_n97_w192, 
            w193=> c0_n97_w193, 
            w194=> c0_n97_w194, 
            w195=> c0_n97_w195, 
            w196=> c0_n97_w196, 
            w197=> c0_n97_w197, 
            w198=> c0_n97_w198, 
            w199=> c0_n97_w199, 
            w200=> c0_n97_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n97_y
   );           
            
neuron_inst_98: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n98_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n98_w1, 
            w2=> c0_n98_w2, 
            w3=> c0_n98_w3, 
            w4=> c0_n98_w4, 
            w5=> c0_n98_w5, 
            w6=> c0_n98_w6, 
            w7=> c0_n98_w7, 
            w8=> c0_n98_w8, 
            w9=> c0_n98_w9, 
            w10=> c0_n98_w10, 
            w11=> c0_n98_w11, 
            w12=> c0_n98_w12, 
            w13=> c0_n98_w13, 
            w14=> c0_n98_w14, 
            w15=> c0_n98_w15, 
            w16=> c0_n98_w16, 
            w17=> c0_n98_w17, 
            w18=> c0_n98_w18, 
            w19=> c0_n98_w19, 
            w20=> c0_n98_w20, 
            w21=> c0_n98_w21, 
            w22=> c0_n98_w22, 
            w23=> c0_n98_w23, 
            w24=> c0_n98_w24, 
            w25=> c0_n98_w25, 
            w26=> c0_n98_w26, 
            w27=> c0_n98_w27, 
            w28=> c0_n98_w28, 
            w29=> c0_n98_w29, 
            w30=> c0_n98_w30, 
            w31=> c0_n98_w31, 
            w32=> c0_n98_w32, 
            w33=> c0_n98_w33, 
            w34=> c0_n98_w34, 
            w35=> c0_n98_w35, 
            w36=> c0_n98_w36, 
            w37=> c0_n98_w37, 
            w38=> c0_n98_w38, 
            w39=> c0_n98_w39, 
            w40=> c0_n98_w40, 
            w41=> c0_n98_w41, 
            w42=> c0_n98_w42, 
            w43=> c0_n98_w43, 
            w44=> c0_n98_w44, 
            w45=> c0_n98_w45, 
            w46=> c0_n98_w46, 
            w47=> c0_n98_w47, 
            w48=> c0_n98_w48, 
            w49=> c0_n98_w49, 
            w50=> c0_n98_w50, 
            w51=> c0_n98_w51, 
            w52=> c0_n98_w52, 
            w53=> c0_n98_w53, 
            w54=> c0_n98_w54, 
            w55=> c0_n98_w55, 
            w56=> c0_n98_w56, 
            w57=> c0_n98_w57, 
            w58=> c0_n98_w58, 
            w59=> c0_n98_w59, 
            w60=> c0_n98_w60, 
            w61=> c0_n98_w61, 
            w62=> c0_n98_w62, 
            w63=> c0_n98_w63, 
            w64=> c0_n98_w64, 
            w65=> c0_n98_w65, 
            w66=> c0_n98_w66, 
            w67=> c0_n98_w67, 
            w68=> c0_n98_w68, 
            w69=> c0_n98_w69, 
            w70=> c0_n98_w70, 
            w71=> c0_n98_w71, 
            w72=> c0_n98_w72, 
            w73=> c0_n98_w73, 
            w74=> c0_n98_w74, 
            w75=> c0_n98_w75, 
            w76=> c0_n98_w76, 
            w77=> c0_n98_w77, 
            w78=> c0_n98_w78, 
            w79=> c0_n98_w79, 
            w80=> c0_n98_w80, 
            w81=> c0_n98_w81, 
            w82=> c0_n98_w82, 
            w83=> c0_n98_w83, 
            w84=> c0_n98_w84, 
            w85=> c0_n98_w85, 
            w86=> c0_n98_w86, 
            w87=> c0_n98_w87, 
            w88=> c0_n98_w88, 
            w89=> c0_n98_w89, 
            w90=> c0_n98_w90, 
            w91=> c0_n98_w91, 
            w92=> c0_n98_w92, 
            w93=> c0_n98_w93, 
            w94=> c0_n98_w94, 
            w95=> c0_n98_w95, 
            w96=> c0_n98_w96, 
            w97=> c0_n98_w97, 
            w98=> c0_n98_w98, 
            w99=> c0_n98_w99, 
            w100=> c0_n98_w100, 
            w101=> c0_n98_w101, 
            w102=> c0_n98_w102, 
            w103=> c0_n98_w103, 
            w104=> c0_n98_w104, 
            w105=> c0_n98_w105, 
            w106=> c0_n98_w106, 
            w107=> c0_n98_w107, 
            w108=> c0_n98_w108, 
            w109=> c0_n98_w109, 
            w110=> c0_n98_w110, 
            w111=> c0_n98_w111, 
            w112=> c0_n98_w112, 
            w113=> c0_n98_w113, 
            w114=> c0_n98_w114, 
            w115=> c0_n98_w115, 
            w116=> c0_n98_w116, 
            w117=> c0_n98_w117, 
            w118=> c0_n98_w118, 
            w119=> c0_n98_w119, 
            w120=> c0_n98_w120, 
            w121=> c0_n98_w121, 
            w122=> c0_n98_w122, 
            w123=> c0_n98_w123, 
            w124=> c0_n98_w124, 
            w125=> c0_n98_w125, 
            w126=> c0_n98_w126, 
            w127=> c0_n98_w127, 
            w128=> c0_n98_w128, 
            w129=> c0_n98_w129, 
            w130=> c0_n98_w130, 
            w131=> c0_n98_w131, 
            w132=> c0_n98_w132, 
            w133=> c0_n98_w133, 
            w134=> c0_n98_w134, 
            w135=> c0_n98_w135, 
            w136=> c0_n98_w136, 
            w137=> c0_n98_w137, 
            w138=> c0_n98_w138, 
            w139=> c0_n98_w139, 
            w140=> c0_n98_w140, 
            w141=> c0_n98_w141, 
            w142=> c0_n98_w142, 
            w143=> c0_n98_w143, 
            w144=> c0_n98_w144, 
            w145=> c0_n98_w145, 
            w146=> c0_n98_w146, 
            w147=> c0_n98_w147, 
            w148=> c0_n98_w148, 
            w149=> c0_n98_w149, 
            w150=> c0_n98_w150, 
            w151=> c0_n98_w151, 
            w152=> c0_n98_w152, 
            w153=> c0_n98_w153, 
            w154=> c0_n98_w154, 
            w155=> c0_n98_w155, 
            w156=> c0_n98_w156, 
            w157=> c0_n98_w157, 
            w158=> c0_n98_w158, 
            w159=> c0_n98_w159, 
            w160=> c0_n98_w160, 
            w161=> c0_n98_w161, 
            w162=> c0_n98_w162, 
            w163=> c0_n98_w163, 
            w164=> c0_n98_w164, 
            w165=> c0_n98_w165, 
            w166=> c0_n98_w166, 
            w167=> c0_n98_w167, 
            w168=> c0_n98_w168, 
            w169=> c0_n98_w169, 
            w170=> c0_n98_w170, 
            w171=> c0_n98_w171, 
            w172=> c0_n98_w172, 
            w173=> c0_n98_w173, 
            w174=> c0_n98_w174, 
            w175=> c0_n98_w175, 
            w176=> c0_n98_w176, 
            w177=> c0_n98_w177, 
            w178=> c0_n98_w178, 
            w179=> c0_n98_w179, 
            w180=> c0_n98_w180, 
            w181=> c0_n98_w181, 
            w182=> c0_n98_w182, 
            w183=> c0_n98_w183, 
            w184=> c0_n98_w184, 
            w185=> c0_n98_w185, 
            w186=> c0_n98_w186, 
            w187=> c0_n98_w187, 
            w188=> c0_n98_w188, 
            w189=> c0_n98_w189, 
            w190=> c0_n98_w190, 
            w191=> c0_n98_w191, 
            w192=> c0_n98_w192, 
            w193=> c0_n98_w193, 
            w194=> c0_n98_w194, 
            w195=> c0_n98_w195, 
            w196=> c0_n98_w196, 
            w197=> c0_n98_w197, 
            w198=> c0_n98_w198, 
            w199=> c0_n98_w199, 
            w200=> c0_n98_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n98_y
   );           
            
neuron_inst_99: ENTITY work.neuron_comb_ReLU_200n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n99_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            x101=> x101, 
            x102=> x102, 
            x103=> x103, 
            x104=> x104, 
            x105=> x105, 
            x106=> x106, 
            x107=> x107, 
            x108=> x108, 
            x109=> x109, 
            x110=> x110, 
            x111=> x111, 
            x112=> x112, 
            x113=> x113, 
            x114=> x114, 
            x115=> x115, 
            x116=> x116, 
            x117=> x117, 
            x118=> x118, 
            x119=> x119, 
            x120=> x120, 
            x121=> x121, 
            x122=> x122, 
            x123=> x123, 
            x124=> x124, 
            x125=> x125, 
            x126=> x126, 
            x127=> x127, 
            x128=> x128, 
            x129=> x129, 
            x130=> x130, 
            x131=> x131, 
            x132=> x132, 
            x133=> x133, 
            x134=> x134, 
            x135=> x135, 
            x136=> x136, 
            x137=> x137, 
            x138=> x138, 
            x139=> x139, 
            x140=> x140, 
            x141=> x141, 
            x142=> x142, 
            x143=> x143, 
            x144=> x144, 
            x145=> x145, 
            x146=> x146, 
            x147=> x147, 
            x148=> x148, 
            x149=> x149, 
            x150=> x150, 
            x151=> x151, 
            x152=> x152, 
            x153=> x153, 
            x154=> x154, 
            x155=> x155, 
            x156=> x156, 
            x157=> x157, 
            x158=> x158, 
            x159=> x159, 
            x160=> x160, 
            x161=> x161, 
            x162=> x162, 
            x163=> x163, 
            x164=> x164, 
            x165=> x165, 
            x166=> x166, 
            x167=> x167, 
            x168=> x168, 
            x169=> x169, 
            x170=> x170, 
            x171=> x171, 
            x172=> x172, 
            x173=> x173, 
            x174=> x174, 
            x175=> x175, 
            x176=> x176, 
            x177=> x177, 
            x178=> x178, 
            x179=> x179, 
            x180=> x180, 
            x181=> x181, 
            x182=> x182, 
            x183=> x183, 
            x184=> x184, 
            x185=> x185, 
            x186=> x186, 
            x187=> x187, 
            x188=> x188, 
            x189=> x189, 
            x190=> x190, 
            x191=> x191, 
            x192=> x192, 
            x193=> x193, 
            x194=> x194, 
            x195=> x195, 
            x196=> x196, 
            x197=> x197, 
            x198=> x198, 
            x199=> x199, 
            x200=> x200, 
            w1=> c0_n99_w1, 
            w2=> c0_n99_w2, 
            w3=> c0_n99_w3, 
            w4=> c0_n99_w4, 
            w5=> c0_n99_w5, 
            w6=> c0_n99_w6, 
            w7=> c0_n99_w7, 
            w8=> c0_n99_w8, 
            w9=> c0_n99_w9, 
            w10=> c0_n99_w10, 
            w11=> c0_n99_w11, 
            w12=> c0_n99_w12, 
            w13=> c0_n99_w13, 
            w14=> c0_n99_w14, 
            w15=> c0_n99_w15, 
            w16=> c0_n99_w16, 
            w17=> c0_n99_w17, 
            w18=> c0_n99_w18, 
            w19=> c0_n99_w19, 
            w20=> c0_n99_w20, 
            w21=> c0_n99_w21, 
            w22=> c0_n99_w22, 
            w23=> c0_n99_w23, 
            w24=> c0_n99_w24, 
            w25=> c0_n99_w25, 
            w26=> c0_n99_w26, 
            w27=> c0_n99_w27, 
            w28=> c0_n99_w28, 
            w29=> c0_n99_w29, 
            w30=> c0_n99_w30, 
            w31=> c0_n99_w31, 
            w32=> c0_n99_w32, 
            w33=> c0_n99_w33, 
            w34=> c0_n99_w34, 
            w35=> c0_n99_w35, 
            w36=> c0_n99_w36, 
            w37=> c0_n99_w37, 
            w38=> c0_n99_w38, 
            w39=> c0_n99_w39, 
            w40=> c0_n99_w40, 
            w41=> c0_n99_w41, 
            w42=> c0_n99_w42, 
            w43=> c0_n99_w43, 
            w44=> c0_n99_w44, 
            w45=> c0_n99_w45, 
            w46=> c0_n99_w46, 
            w47=> c0_n99_w47, 
            w48=> c0_n99_w48, 
            w49=> c0_n99_w49, 
            w50=> c0_n99_w50, 
            w51=> c0_n99_w51, 
            w52=> c0_n99_w52, 
            w53=> c0_n99_w53, 
            w54=> c0_n99_w54, 
            w55=> c0_n99_w55, 
            w56=> c0_n99_w56, 
            w57=> c0_n99_w57, 
            w58=> c0_n99_w58, 
            w59=> c0_n99_w59, 
            w60=> c0_n99_w60, 
            w61=> c0_n99_w61, 
            w62=> c0_n99_w62, 
            w63=> c0_n99_w63, 
            w64=> c0_n99_w64, 
            w65=> c0_n99_w65, 
            w66=> c0_n99_w66, 
            w67=> c0_n99_w67, 
            w68=> c0_n99_w68, 
            w69=> c0_n99_w69, 
            w70=> c0_n99_w70, 
            w71=> c0_n99_w71, 
            w72=> c0_n99_w72, 
            w73=> c0_n99_w73, 
            w74=> c0_n99_w74, 
            w75=> c0_n99_w75, 
            w76=> c0_n99_w76, 
            w77=> c0_n99_w77, 
            w78=> c0_n99_w78, 
            w79=> c0_n99_w79, 
            w80=> c0_n99_w80, 
            w81=> c0_n99_w81, 
            w82=> c0_n99_w82, 
            w83=> c0_n99_w83, 
            w84=> c0_n99_w84, 
            w85=> c0_n99_w85, 
            w86=> c0_n99_w86, 
            w87=> c0_n99_w87, 
            w88=> c0_n99_w88, 
            w89=> c0_n99_w89, 
            w90=> c0_n99_w90, 
            w91=> c0_n99_w91, 
            w92=> c0_n99_w92, 
            w93=> c0_n99_w93, 
            w94=> c0_n99_w94, 
            w95=> c0_n99_w95, 
            w96=> c0_n99_w96, 
            w97=> c0_n99_w97, 
            w98=> c0_n99_w98, 
            w99=> c0_n99_w99, 
            w100=> c0_n99_w100, 
            w101=> c0_n99_w101, 
            w102=> c0_n99_w102, 
            w103=> c0_n99_w103, 
            w104=> c0_n99_w104, 
            w105=> c0_n99_w105, 
            w106=> c0_n99_w106, 
            w107=> c0_n99_w107, 
            w108=> c0_n99_w108, 
            w109=> c0_n99_w109, 
            w110=> c0_n99_w110, 
            w111=> c0_n99_w111, 
            w112=> c0_n99_w112, 
            w113=> c0_n99_w113, 
            w114=> c0_n99_w114, 
            w115=> c0_n99_w115, 
            w116=> c0_n99_w116, 
            w117=> c0_n99_w117, 
            w118=> c0_n99_w118, 
            w119=> c0_n99_w119, 
            w120=> c0_n99_w120, 
            w121=> c0_n99_w121, 
            w122=> c0_n99_w122, 
            w123=> c0_n99_w123, 
            w124=> c0_n99_w124, 
            w125=> c0_n99_w125, 
            w126=> c0_n99_w126, 
            w127=> c0_n99_w127, 
            w128=> c0_n99_w128, 
            w129=> c0_n99_w129, 
            w130=> c0_n99_w130, 
            w131=> c0_n99_w131, 
            w132=> c0_n99_w132, 
            w133=> c0_n99_w133, 
            w134=> c0_n99_w134, 
            w135=> c0_n99_w135, 
            w136=> c0_n99_w136, 
            w137=> c0_n99_w137, 
            w138=> c0_n99_w138, 
            w139=> c0_n99_w139, 
            w140=> c0_n99_w140, 
            w141=> c0_n99_w141, 
            w142=> c0_n99_w142, 
            w143=> c0_n99_w143, 
            w144=> c0_n99_w144, 
            w145=> c0_n99_w145, 
            w146=> c0_n99_w146, 
            w147=> c0_n99_w147, 
            w148=> c0_n99_w148, 
            w149=> c0_n99_w149, 
            w150=> c0_n99_w150, 
            w151=> c0_n99_w151, 
            w152=> c0_n99_w152, 
            w153=> c0_n99_w153, 
            w154=> c0_n99_w154, 
            w155=> c0_n99_w155, 
            w156=> c0_n99_w156, 
            w157=> c0_n99_w157, 
            w158=> c0_n99_w158, 
            w159=> c0_n99_w159, 
            w160=> c0_n99_w160, 
            w161=> c0_n99_w161, 
            w162=> c0_n99_w162, 
            w163=> c0_n99_w163, 
            w164=> c0_n99_w164, 
            w165=> c0_n99_w165, 
            w166=> c0_n99_w166, 
            w167=> c0_n99_w167, 
            w168=> c0_n99_w168, 
            w169=> c0_n99_w169, 
            w170=> c0_n99_w170, 
            w171=> c0_n99_w171, 
            w172=> c0_n99_w172, 
            w173=> c0_n99_w173, 
            w174=> c0_n99_w174, 
            w175=> c0_n99_w175, 
            w176=> c0_n99_w176, 
            w177=> c0_n99_w177, 
            w178=> c0_n99_w178, 
            w179=> c0_n99_w179, 
            w180=> c0_n99_w180, 
            w181=> c0_n99_w181, 
            w182=> c0_n99_w182, 
            w183=> c0_n99_w183, 
            w184=> c0_n99_w184, 
            w185=> c0_n99_w185, 
            w186=> c0_n99_w186, 
            w187=> c0_n99_w187, 
            w188=> c0_n99_w188, 
            w189=> c0_n99_w189, 
            w190=> c0_n99_w190, 
            w191=> c0_n99_w191, 
            w192=> c0_n99_w192, 
            w193=> c0_n99_w193, 
            w194=> c0_n99_w194, 
            w195=> c0_n99_w195, 
            w196=> c0_n99_w196, 
            w197=> c0_n99_w197, 
            w198=> c0_n99_w198, 
            w199=> c0_n99_w199, 
            w200=> c0_n99_w200, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n99_y
   );           
             
END ARCHITECTURE;
