LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada3_Sigmoid_5neuron_8bits_30n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c3_n0_bias, c3_n1_bias, c3_n2_bias, c3_n3_bias, c3_n4_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, c3_n0_w1, c3_n0_w2, c3_n0_w3, c3_n0_w4, c3_n0_w5, c3_n0_w6, c3_n0_w7, c3_n0_w8, c3_n0_w9, c3_n0_w10, c3_n0_w11, c3_n0_w12, c3_n0_w13, c3_n0_w14, c3_n0_w15, c3_n0_w16, c3_n0_w17, c3_n0_w18, c3_n0_w19, c3_n0_w20, c3_n0_w21, c3_n0_w22, c3_n0_w23, c3_n0_w24, c3_n0_w25, c3_n0_w26, c3_n0_w27, c3_n0_w28, c3_n0_w29, c3_n0_w30, c3_n1_w1, c3_n1_w2, c3_n1_w3, c3_n1_w4, c3_n1_w5, c3_n1_w6, c3_n1_w7, c3_n1_w8, c3_n1_w9, c3_n1_w10, c3_n1_w11, c3_n1_w12, c3_n1_w13, c3_n1_w14, c3_n1_w15, c3_n1_w16, c3_n1_w17, c3_n1_w18, c3_n1_w19, c3_n1_w20, c3_n1_w21, c3_n1_w22, c3_n1_w23, c3_n1_w24, c3_n1_w25, c3_n1_w26, c3_n1_w27, c3_n1_w28, c3_n1_w29, c3_n1_w30, c3_n2_w1, c3_n2_w2, c3_n2_w3, c3_n2_w4, c3_n2_w5, c3_n2_w6, c3_n2_w7, c3_n2_w8, c3_n2_w9, c3_n2_w10, c3_n2_w11, c3_n2_w12, c3_n2_w13, c3_n2_w14, c3_n2_w15, c3_n2_w16, c3_n2_w17, c3_n2_w18, c3_n2_w19, c3_n2_w20, c3_n2_w21, c3_n2_w22, c3_n2_w23, c3_n2_w24, c3_n2_w25, c3_n2_w26, c3_n2_w27, c3_n2_w28, c3_n2_w29, c3_n2_w30, c3_n3_w1, c3_n3_w2, c3_n3_w3, c3_n3_w4, c3_n3_w5, c3_n3_w6, c3_n3_w7, c3_n3_w8, c3_n3_w9, c3_n3_w10, c3_n3_w11, c3_n3_w12, c3_n3_w13, c3_n3_w14, c3_n3_w15, c3_n3_w16, c3_n3_w17, c3_n3_w18, c3_n3_w19, c3_n3_w20, c3_n3_w21, c3_n3_w22, c3_n3_w23, c3_n3_w24, c3_n3_w25, c3_n3_w26, c3_n3_w27, c3_n3_w28, c3_n3_w29, c3_n3_w30, c3_n4_w1, c3_n4_w2, c3_n4_w3, c3_n4_w4, c3_n4_w5, c3_n4_w6, c3_n4_w7, c3_n4_w8, c3_n4_w9, c3_n4_w10, c3_n4_w11, c3_n4_w12, c3_n4_w13, c3_n4_w14, c3_n4_w15, c3_n4_w16, c3_n4_w17, c3_n4_w18, c3_n4_w19, c3_n4_w20, c3_n4_w21, c3_n4_w22, c3_n4_w23, c3_n4_w24, c3_n4_w25, c3_n4_w26, c3_n4_w27, c3_n4_w28, c3_n4_w29, c3_n4_w30: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c3_n0_y, c3_n1_y, c3_n2_y, c3_n3_y, c3_n4_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada3_Sigmoid_5neuron_8bits_30n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_Sigmoid_30n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c3_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            w1=> c3_n0_w1, 
            w2=> c3_n0_w2, 
            w3=> c3_n0_w3, 
            w4=> c3_n0_w4, 
            w5=> c3_n0_w5, 
            w6=> c3_n0_w6, 
            w7=> c3_n0_w7, 
            w8=> c3_n0_w8, 
            w9=> c3_n0_w9, 
            w10=> c3_n0_w10, 
            w11=> c3_n0_w11, 
            w12=> c3_n0_w12, 
            w13=> c3_n0_w13, 
            w14=> c3_n0_w14, 
            w15=> c3_n0_w15, 
            w16=> c3_n0_w16, 
            w17=> c3_n0_w17, 
            w18=> c3_n0_w18, 
            w19=> c3_n0_w19, 
            w20=> c3_n0_w20, 
            w21=> c3_n0_w21, 
            w22=> c3_n0_w22, 
            w23=> c3_n0_w23, 
            w24=> c3_n0_w24, 
            w25=> c3_n0_w25, 
            w26=> c3_n0_w26, 
            w27=> c3_n0_w27, 
            w28=> c3_n0_w28, 
            w29=> c3_n0_w29, 
            w30=> c3_n0_w30, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c3_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_Sigmoid_30n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c3_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            w1=> c3_n1_w1, 
            w2=> c3_n1_w2, 
            w3=> c3_n1_w3, 
            w4=> c3_n1_w4, 
            w5=> c3_n1_w5, 
            w6=> c3_n1_w6, 
            w7=> c3_n1_w7, 
            w8=> c3_n1_w8, 
            w9=> c3_n1_w9, 
            w10=> c3_n1_w10, 
            w11=> c3_n1_w11, 
            w12=> c3_n1_w12, 
            w13=> c3_n1_w13, 
            w14=> c3_n1_w14, 
            w15=> c3_n1_w15, 
            w16=> c3_n1_w16, 
            w17=> c3_n1_w17, 
            w18=> c3_n1_w18, 
            w19=> c3_n1_w19, 
            w20=> c3_n1_w20, 
            w21=> c3_n1_w21, 
            w22=> c3_n1_w22, 
            w23=> c3_n1_w23, 
            w24=> c3_n1_w24, 
            w25=> c3_n1_w25, 
            w26=> c3_n1_w26, 
            w27=> c3_n1_w27, 
            w28=> c3_n1_w28, 
            w29=> c3_n1_w29, 
            w30=> c3_n1_w30, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c3_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_Sigmoid_30n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c3_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            w1=> c3_n2_w1, 
            w2=> c3_n2_w2, 
            w3=> c3_n2_w3, 
            w4=> c3_n2_w4, 
            w5=> c3_n2_w5, 
            w6=> c3_n2_w6, 
            w7=> c3_n2_w7, 
            w8=> c3_n2_w8, 
            w9=> c3_n2_w9, 
            w10=> c3_n2_w10, 
            w11=> c3_n2_w11, 
            w12=> c3_n2_w12, 
            w13=> c3_n2_w13, 
            w14=> c3_n2_w14, 
            w15=> c3_n2_w15, 
            w16=> c3_n2_w16, 
            w17=> c3_n2_w17, 
            w18=> c3_n2_w18, 
            w19=> c3_n2_w19, 
            w20=> c3_n2_w20, 
            w21=> c3_n2_w21, 
            w22=> c3_n2_w22, 
            w23=> c3_n2_w23, 
            w24=> c3_n2_w24, 
            w25=> c3_n2_w25, 
            w26=> c3_n2_w26, 
            w27=> c3_n2_w27, 
            w28=> c3_n2_w28, 
            w29=> c3_n2_w29, 
            w30=> c3_n2_w30, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c3_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_Sigmoid_30n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c3_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            w1=> c3_n3_w1, 
            w2=> c3_n3_w2, 
            w3=> c3_n3_w3, 
            w4=> c3_n3_w4, 
            w5=> c3_n3_w5, 
            w6=> c3_n3_w6, 
            w7=> c3_n3_w7, 
            w8=> c3_n3_w8, 
            w9=> c3_n3_w9, 
            w10=> c3_n3_w10, 
            w11=> c3_n3_w11, 
            w12=> c3_n3_w12, 
            w13=> c3_n3_w13, 
            w14=> c3_n3_w14, 
            w15=> c3_n3_w15, 
            w16=> c3_n3_w16, 
            w17=> c3_n3_w17, 
            w18=> c3_n3_w18, 
            w19=> c3_n3_w19, 
            w20=> c3_n3_w20, 
            w21=> c3_n3_w21, 
            w22=> c3_n3_w22, 
            w23=> c3_n3_w23, 
            w24=> c3_n3_w24, 
            w25=> c3_n3_w25, 
            w26=> c3_n3_w26, 
            w27=> c3_n3_w27, 
            w28=> c3_n3_w28, 
            w29=> c3_n3_w29, 
            w30=> c3_n3_w30, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c3_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_Sigmoid_30n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c3_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            w1=> c3_n4_w1, 
            w2=> c3_n4_w2, 
            w3=> c3_n4_w3, 
            w4=> c3_n4_w4, 
            w5=> c3_n4_w5, 
            w6=> c3_n4_w6, 
            w7=> c3_n4_w7, 
            w8=> c3_n4_w8, 
            w9=> c3_n4_w9, 
            w10=> c3_n4_w10, 
            w11=> c3_n4_w11, 
            w12=> c3_n4_w12, 
            w13=> c3_n4_w13, 
            w14=> c3_n4_w14, 
            w15=> c3_n4_w15, 
            w16=> c3_n4_w16, 
            w17=> c3_n4_w17, 
            w18=> c3_n4_w18, 
            w19=> c3_n4_w19, 
            w20=> c3_n4_w20, 
            w21=> c3_n4_w21, 
            w22=> c3_n4_w22, 
            w23=> c3_n4_w23, 
            w24=> c3_n4_w24, 
            w25=> c3_n4_w25, 
            w26=> c3_n4_w26, 
            w27=> c3_n4_w27, 
            w28=> c3_n4_w28, 
            w29=> c3_n4_w29, 
            w30=> c3_n4_w30, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c3_n4_y
   );           
             
END ARCHITECTURE;
