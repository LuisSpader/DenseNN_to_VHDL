LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada0_ReLU_15neuron_8bits_64n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c0_n0_bias, c0_n1_bias, c0_n2_bias, c0_n3_bias, c0_n4_bias, c0_n5_bias, c0_n6_bias, c0_n7_bias, c0_n8_bias, c0_n9_bias, c0_n10_bias, c0_n11_bias, c0_n12_bias, c0_n13_bias, c0_n14_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, c0_n0_w1, c0_n0_w2, c0_n0_w3, c0_n0_w4, c0_n0_w5, c0_n0_w6, c0_n0_w7, c0_n0_w8, c0_n0_w9, c0_n0_w10, c0_n0_w11, c0_n0_w12, c0_n0_w13, c0_n0_w14, c0_n0_w15, c0_n0_w16, c0_n0_w17, c0_n0_w18, c0_n0_w19, c0_n0_w20, c0_n0_w21, c0_n0_w22, c0_n0_w23, c0_n0_w24, c0_n0_w25, c0_n0_w26, c0_n0_w27, c0_n0_w28, c0_n0_w29, c0_n0_w30, c0_n0_w31, c0_n0_w32, c0_n0_w33, c0_n0_w34, c0_n0_w35, c0_n0_w36, c0_n0_w37, c0_n0_w38, c0_n0_w39, c0_n0_w40, c0_n0_w41, c0_n0_w42, c0_n0_w43, c0_n0_w44, c0_n0_w45, c0_n0_w46, c0_n0_w47, c0_n0_w48, c0_n0_w49, c0_n0_w50, c0_n0_w51, c0_n0_w52, c0_n0_w53, c0_n0_w54, c0_n0_w55, c0_n0_w56, c0_n0_w57, c0_n0_w58, c0_n0_w59, c0_n0_w60, c0_n0_w61, c0_n0_w62, c0_n0_w63, c0_n0_w64, c0_n1_w1, c0_n1_w2, c0_n1_w3, c0_n1_w4, c0_n1_w5, c0_n1_w6, c0_n1_w7, c0_n1_w8, c0_n1_w9, c0_n1_w10, c0_n1_w11, c0_n1_w12, c0_n1_w13, c0_n1_w14, c0_n1_w15, c0_n1_w16, c0_n1_w17, c0_n1_w18, c0_n1_w19, c0_n1_w20, c0_n1_w21, c0_n1_w22, c0_n1_w23, c0_n1_w24, c0_n1_w25, c0_n1_w26, c0_n1_w27, c0_n1_w28, c0_n1_w29, c0_n1_w30, c0_n1_w31, c0_n1_w32, c0_n1_w33, c0_n1_w34, c0_n1_w35, c0_n1_w36, c0_n1_w37, c0_n1_w38, c0_n1_w39, c0_n1_w40, c0_n1_w41, c0_n1_w42, c0_n1_w43, c0_n1_w44, c0_n1_w45, c0_n1_w46, c0_n1_w47, c0_n1_w48, c0_n1_w49, c0_n1_w50, c0_n1_w51, c0_n1_w52, c0_n1_w53, c0_n1_w54, c0_n1_w55, c0_n1_w56, c0_n1_w57, c0_n1_w58, c0_n1_w59, c0_n1_w60, c0_n1_w61, c0_n1_w62, c0_n1_w63, c0_n1_w64, c0_n2_w1, c0_n2_w2, c0_n2_w3, c0_n2_w4, c0_n2_w5, c0_n2_w6, c0_n2_w7, c0_n2_w8, c0_n2_w9, c0_n2_w10, c0_n2_w11, c0_n2_w12, c0_n2_w13, c0_n2_w14, c0_n2_w15, c0_n2_w16, c0_n2_w17, c0_n2_w18, c0_n2_w19, c0_n2_w20, c0_n2_w21, c0_n2_w22, c0_n2_w23, c0_n2_w24, c0_n2_w25, c0_n2_w26, c0_n2_w27, c0_n2_w28, c0_n2_w29, c0_n2_w30, c0_n2_w31, c0_n2_w32, c0_n2_w33, c0_n2_w34, c0_n2_w35, c0_n2_w36, c0_n2_w37, c0_n2_w38, c0_n2_w39, c0_n2_w40, c0_n2_w41, c0_n2_w42, c0_n2_w43, c0_n2_w44, c0_n2_w45, c0_n2_w46, c0_n2_w47, c0_n2_w48, c0_n2_w49, c0_n2_w50, c0_n2_w51, c0_n2_w52, c0_n2_w53, c0_n2_w54, c0_n2_w55, c0_n2_w56, c0_n2_w57, c0_n2_w58, c0_n2_w59, c0_n2_w60, c0_n2_w61, c0_n2_w62, c0_n2_w63, c0_n2_w64, c0_n3_w1, c0_n3_w2, c0_n3_w3, c0_n3_w4, c0_n3_w5, c0_n3_w6, c0_n3_w7, c0_n3_w8, c0_n3_w9, c0_n3_w10, c0_n3_w11, c0_n3_w12, c0_n3_w13, c0_n3_w14, c0_n3_w15, c0_n3_w16, c0_n3_w17, c0_n3_w18, c0_n3_w19, c0_n3_w20, c0_n3_w21, c0_n3_w22, c0_n3_w23, c0_n3_w24, c0_n3_w25, c0_n3_w26, c0_n3_w27, c0_n3_w28, c0_n3_w29, c0_n3_w30, c0_n3_w31, c0_n3_w32, c0_n3_w33, c0_n3_w34, c0_n3_w35, c0_n3_w36, c0_n3_w37, c0_n3_w38, c0_n3_w39, c0_n3_w40, c0_n3_w41, c0_n3_w42, c0_n3_w43, c0_n3_w44, c0_n3_w45, c0_n3_w46, c0_n3_w47, c0_n3_w48, c0_n3_w49, c0_n3_w50, c0_n3_w51, c0_n3_w52, c0_n3_w53, c0_n3_w54, c0_n3_w55, c0_n3_w56, c0_n3_w57, c0_n3_w58, c0_n3_w59, c0_n3_w60, c0_n3_w61, c0_n3_w62, c0_n3_w63, c0_n3_w64, c0_n4_w1, c0_n4_w2, c0_n4_w3, c0_n4_w4, c0_n4_w5, c0_n4_w6, c0_n4_w7, c0_n4_w8, c0_n4_w9, c0_n4_w10, c0_n4_w11, c0_n4_w12, c0_n4_w13, c0_n4_w14, c0_n4_w15, c0_n4_w16, c0_n4_w17, c0_n4_w18, c0_n4_w19, c0_n4_w20, c0_n4_w21, c0_n4_w22, c0_n4_w23, c0_n4_w24, c0_n4_w25, c0_n4_w26, c0_n4_w27, c0_n4_w28, c0_n4_w29, c0_n4_w30, c0_n4_w31, c0_n4_w32, c0_n4_w33, c0_n4_w34, c0_n4_w35, c0_n4_w36, c0_n4_w37, c0_n4_w38, c0_n4_w39, c0_n4_w40, c0_n4_w41, c0_n4_w42, c0_n4_w43, c0_n4_w44, c0_n4_w45, c0_n4_w46, c0_n4_w47, c0_n4_w48, c0_n4_w49, c0_n4_w50, c0_n4_w51, c0_n4_w52, c0_n4_w53, c0_n4_w54, c0_n4_w55, c0_n4_w56, c0_n4_w57, c0_n4_w58, c0_n4_w59, c0_n4_w60, c0_n4_w61, c0_n4_w62, c0_n4_w63, c0_n4_w64, c0_n5_w1, c0_n5_w2, c0_n5_w3, c0_n5_w4, c0_n5_w5, c0_n5_w6, c0_n5_w7, c0_n5_w8, c0_n5_w9, c0_n5_w10, c0_n5_w11, c0_n5_w12, c0_n5_w13, c0_n5_w14, c0_n5_w15, c0_n5_w16, c0_n5_w17, c0_n5_w18, c0_n5_w19, c0_n5_w20, c0_n5_w21, c0_n5_w22, c0_n5_w23, c0_n5_w24, c0_n5_w25, c0_n5_w26, c0_n5_w27, c0_n5_w28, c0_n5_w29, c0_n5_w30, c0_n5_w31, c0_n5_w32, c0_n5_w33, c0_n5_w34, c0_n5_w35, c0_n5_w36, c0_n5_w37, c0_n5_w38, c0_n5_w39, c0_n5_w40, c0_n5_w41, c0_n5_w42, c0_n5_w43, c0_n5_w44, c0_n5_w45, c0_n5_w46, c0_n5_w47, c0_n5_w48, c0_n5_w49, c0_n5_w50, c0_n5_w51, c0_n5_w52, c0_n5_w53, c0_n5_w54, c0_n5_w55, c0_n5_w56, c0_n5_w57, c0_n5_w58, c0_n5_w59, c0_n5_w60, c0_n5_w61, c0_n5_w62, c0_n5_w63, c0_n5_w64, c0_n6_w1, c0_n6_w2, c0_n6_w3, c0_n6_w4, c0_n6_w5, c0_n6_w6, c0_n6_w7, c0_n6_w8, c0_n6_w9, c0_n6_w10, c0_n6_w11, c0_n6_w12, c0_n6_w13, c0_n6_w14, c0_n6_w15, c0_n6_w16, c0_n6_w17, c0_n6_w18, c0_n6_w19, c0_n6_w20, c0_n6_w21, c0_n6_w22, c0_n6_w23, c0_n6_w24, c0_n6_w25, c0_n6_w26, c0_n6_w27, c0_n6_w28, c0_n6_w29, c0_n6_w30, c0_n6_w31, c0_n6_w32, c0_n6_w33, c0_n6_w34, c0_n6_w35, c0_n6_w36, c0_n6_w37, c0_n6_w38, c0_n6_w39, c0_n6_w40, c0_n6_w41, c0_n6_w42, c0_n6_w43, c0_n6_w44, c0_n6_w45, c0_n6_w46, c0_n6_w47, c0_n6_w48, c0_n6_w49, c0_n6_w50, c0_n6_w51, c0_n6_w52, c0_n6_w53, c0_n6_w54, c0_n6_w55, c0_n6_w56, c0_n6_w57, c0_n6_w58, c0_n6_w59, c0_n6_w60, c0_n6_w61, c0_n6_w62, c0_n6_w63, c0_n6_w64, c0_n7_w1, c0_n7_w2, c0_n7_w3, c0_n7_w4, c0_n7_w5, c0_n7_w6, c0_n7_w7, c0_n7_w8, c0_n7_w9, c0_n7_w10, c0_n7_w11, c0_n7_w12, c0_n7_w13, c0_n7_w14, c0_n7_w15, c0_n7_w16, c0_n7_w17, c0_n7_w18, c0_n7_w19, c0_n7_w20, c0_n7_w21, c0_n7_w22, c0_n7_w23, c0_n7_w24, c0_n7_w25, c0_n7_w26, c0_n7_w27, c0_n7_w28, c0_n7_w29, c0_n7_w30, c0_n7_w31, c0_n7_w32, c0_n7_w33, c0_n7_w34, c0_n7_w35, c0_n7_w36, c0_n7_w37, c0_n7_w38, c0_n7_w39, c0_n7_w40, c0_n7_w41, c0_n7_w42, c0_n7_w43, c0_n7_w44, c0_n7_w45, c0_n7_w46, c0_n7_w47, c0_n7_w48, c0_n7_w49, c0_n7_w50, c0_n7_w51, c0_n7_w52, c0_n7_w53, c0_n7_w54, c0_n7_w55, c0_n7_w56, c0_n7_w57, c0_n7_w58, c0_n7_w59, c0_n7_w60, c0_n7_w61, c0_n7_w62, c0_n7_w63, c0_n7_w64, c0_n8_w1, c0_n8_w2, c0_n8_w3, c0_n8_w4, c0_n8_w5, c0_n8_w6, c0_n8_w7, c0_n8_w8, c0_n8_w9, c0_n8_w10, c0_n8_w11, c0_n8_w12, c0_n8_w13, c0_n8_w14, c0_n8_w15, c0_n8_w16, c0_n8_w17, c0_n8_w18, c0_n8_w19, c0_n8_w20, c0_n8_w21, c0_n8_w22, c0_n8_w23, c0_n8_w24, c0_n8_w25, c0_n8_w26, c0_n8_w27, c0_n8_w28, c0_n8_w29, c0_n8_w30, c0_n8_w31, c0_n8_w32, c0_n8_w33, c0_n8_w34, c0_n8_w35, c0_n8_w36, c0_n8_w37, c0_n8_w38, c0_n8_w39, c0_n8_w40, c0_n8_w41, c0_n8_w42, c0_n8_w43, c0_n8_w44, c0_n8_w45, c0_n8_w46, c0_n8_w47, c0_n8_w48, c0_n8_w49, c0_n8_w50, c0_n8_w51, c0_n8_w52, c0_n8_w53, c0_n8_w54, c0_n8_w55, c0_n8_w56, c0_n8_w57, c0_n8_w58, c0_n8_w59, c0_n8_w60, c0_n8_w61, c0_n8_w62, c0_n8_w63, c0_n8_w64, c0_n9_w1, c0_n9_w2, c0_n9_w3, c0_n9_w4, c0_n9_w5, c0_n9_w6, c0_n9_w7, c0_n9_w8, c0_n9_w9, c0_n9_w10, c0_n9_w11, c0_n9_w12, c0_n9_w13, c0_n9_w14, c0_n9_w15, c0_n9_w16, c0_n9_w17, c0_n9_w18, c0_n9_w19, c0_n9_w20, c0_n9_w21, c0_n9_w22, c0_n9_w23, c0_n9_w24, c0_n9_w25, c0_n9_w26, c0_n9_w27, c0_n9_w28, c0_n9_w29, c0_n9_w30, c0_n9_w31, c0_n9_w32, c0_n9_w33, c0_n9_w34, c0_n9_w35, c0_n9_w36, c0_n9_w37, c0_n9_w38, c0_n9_w39, c0_n9_w40, c0_n9_w41, c0_n9_w42, c0_n9_w43, c0_n9_w44, c0_n9_w45, c0_n9_w46, c0_n9_w47, c0_n9_w48, c0_n9_w49, c0_n9_w50, c0_n9_w51, c0_n9_w52, c0_n9_w53, c0_n9_w54, c0_n9_w55, c0_n9_w56, c0_n9_w57, c0_n9_w58, c0_n9_w59, c0_n9_w60, c0_n9_w61, c0_n9_w62, c0_n9_w63, c0_n9_w64, c0_n10_w1, c0_n10_w2, c0_n10_w3, c0_n10_w4, c0_n10_w5, c0_n10_w6, c0_n10_w7, c0_n10_w8, c0_n10_w9, c0_n10_w10, c0_n10_w11, c0_n10_w12, c0_n10_w13, c0_n10_w14, c0_n10_w15, c0_n10_w16, c0_n10_w17, c0_n10_w18, c0_n10_w19, c0_n10_w20, c0_n10_w21, c0_n10_w22, c0_n10_w23, c0_n10_w24, c0_n10_w25, c0_n10_w26, c0_n10_w27, c0_n10_w28, c0_n10_w29, c0_n10_w30, c0_n10_w31, c0_n10_w32, c0_n10_w33, c0_n10_w34, c0_n10_w35, c0_n10_w36, c0_n10_w37, c0_n10_w38, c0_n10_w39, c0_n10_w40, c0_n10_w41, c0_n10_w42, c0_n10_w43, c0_n10_w44, c0_n10_w45, c0_n10_w46, c0_n10_w47, c0_n10_w48, c0_n10_w49, c0_n10_w50, c0_n10_w51, c0_n10_w52, c0_n10_w53, c0_n10_w54, c0_n10_w55, c0_n10_w56, c0_n10_w57, c0_n10_w58, c0_n10_w59, c0_n10_w60, c0_n10_w61, c0_n10_w62, c0_n10_w63, c0_n10_w64, c0_n11_w1, c0_n11_w2, c0_n11_w3, c0_n11_w4, c0_n11_w5, c0_n11_w6, c0_n11_w7, c0_n11_w8, c0_n11_w9, c0_n11_w10, c0_n11_w11, c0_n11_w12, c0_n11_w13, c0_n11_w14, c0_n11_w15, c0_n11_w16, c0_n11_w17, c0_n11_w18, c0_n11_w19, c0_n11_w20, c0_n11_w21, c0_n11_w22, c0_n11_w23, c0_n11_w24, c0_n11_w25, c0_n11_w26, c0_n11_w27, c0_n11_w28, c0_n11_w29, c0_n11_w30, c0_n11_w31, c0_n11_w32, c0_n11_w33, c0_n11_w34, c0_n11_w35, c0_n11_w36, c0_n11_w37, c0_n11_w38, c0_n11_w39, c0_n11_w40, c0_n11_w41, c0_n11_w42, c0_n11_w43, c0_n11_w44, c0_n11_w45, c0_n11_w46, c0_n11_w47, c0_n11_w48, c0_n11_w49, c0_n11_w50, c0_n11_w51, c0_n11_w52, c0_n11_w53, c0_n11_w54, c0_n11_w55, c0_n11_w56, c0_n11_w57, c0_n11_w58, c0_n11_w59, c0_n11_w60, c0_n11_w61, c0_n11_w62, c0_n11_w63, c0_n11_w64, c0_n12_w1, c0_n12_w2, c0_n12_w3, c0_n12_w4, c0_n12_w5, c0_n12_w6, c0_n12_w7, c0_n12_w8, c0_n12_w9, c0_n12_w10, c0_n12_w11, c0_n12_w12, c0_n12_w13, c0_n12_w14, c0_n12_w15, c0_n12_w16, c0_n12_w17, c0_n12_w18, c0_n12_w19, c0_n12_w20, c0_n12_w21, c0_n12_w22, c0_n12_w23, c0_n12_w24, c0_n12_w25, c0_n12_w26, c0_n12_w27, c0_n12_w28, c0_n12_w29, c0_n12_w30, c0_n12_w31, c0_n12_w32, c0_n12_w33, c0_n12_w34, c0_n12_w35, c0_n12_w36, c0_n12_w37, c0_n12_w38, c0_n12_w39, c0_n12_w40, c0_n12_w41, c0_n12_w42, c0_n12_w43, c0_n12_w44, c0_n12_w45, c0_n12_w46, c0_n12_w47, c0_n12_w48, c0_n12_w49, c0_n12_w50, c0_n12_w51, c0_n12_w52, c0_n12_w53, c0_n12_w54, c0_n12_w55, c0_n12_w56, c0_n12_w57, c0_n12_w58, c0_n12_w59, c0_n12_w60, c0_n12_w61, c0_n12_w62, c0_n12_w63, c0_n12_w64, c0_n13_w1, c0_n13_w2, c0_n13_w3, c0_n13_w4, c0_n13_w5, c0_n13_w6, c0_n13_w7, c0_n13_w8, c0_n13_w9, c0_n13_w10, c0_n13_w11, c0_n13_w12, c0_n13_w13, c0_n13_w14, c0_n13_w15, c0_n13_w16, c0_n13_w17, c0_n13_w18, c0_n13_w19, c0_n13_w20, c0_n13_w21, c0_n13_w22, c0_n13_w23, c0_n13_w24, c0_n13_w25, c0_n13_w26, c0_n13_w27, c0_n13_w28, c0_n13_w29, c0_n13_w30, c0_n13_w31, c0_n13_w32, c0_n13_w33, c0_n13_w34, c0_n13_w35, c0_n13_w36, c0_n13_w37, c0_n13_w38, c0_n13_w39, c0_n13_w40, c0_n13_w41, c0_n13_w42, c0_n13_w43, c0_n13_w44, c0_n13_w45, c0_n13_w46, c0_n13_w47, c0_n13_w48, c0_n13_w49, c0_n13_w50, c0_n13_w51, c0_n13_w52, c0_n13_w53, c0_n13_w54, c0_n13_w55, c0_n13_w56, c0_n13_w57, c0_n13_w58, c0_n13_w59, c0_n13_w60, c0_n13_w61, c0_n13_w62, c0_n13_w63, c0_n13_w64, c0_n14_w1, c0_n14_w2, c0_n14_w3, c0_n14_w4, c0_n14_w5, c0_n14_w6, c0_n14_w7, c0_n14_w8, c0_n14_w9, c0_n14_w10, c0_n14_w11, c0_n14_w12, c0_n14_w13, c0_n14_w14, c0_n14_w15, c0_n14_w16, c0_n14_w17, c0_n14_w18, c0_n14_w19, c0_n14_w20, c0_n14_w21, c0_n14_w22, c0_n14_w23, c0_n14_w24, c0_n14_w25, c0_n14_w26, c0_n14_w27, c0_n14_w28, c0_n14_w29, c0_n14_w30, c0_n14_w31, c0_n14_w32, c0_n14_w33, c0_n14_w34, c0_n14_w35, c0_n14_w36, c0_n14_w37, c0_n14_w38, c0_n14_w39, c0_n14_w40, c0_n14_w41, c0_n14_w42, c0_n14_w43, c0_n14_w44, c0_n14_w45, c0_n14_w46, c0_n14_w47, c0_n14_w48, c0_n14_w49, c0_n14_w50, c0_n14_w51, c0_n14_w52, c0_n14_w53, c0_n14_w54, c0_n14_w55, c0_n14_w56, c0_n14_w57, c0_n14_w58, c0_n14_w59, c0_n14_w60, c0_n14_w61, c0_n14_w62, c0_n14_w63, c0_n14_w64: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c0_n0_y, c0_n1_y, c0_n2_y, c0_n3_y, c0_n4_y, c0_n5_y, c0_n6_y, c0_n7_y, c0_n8_y, c0_n9_y, c0_n10_y, c0_n11_y, c0_n12_y, c0_n13_y, c0_n14_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada0_ReLU_15neuron_8bits_64n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n0_w1, 
            w2=> c0_n0_w2, 
            w3=> c0_n0_w3, 
            w4=> c0_n0_w4, 
            w5=> c0_n0_w5, 
            w6=> c0_n0_w6, 
            w7=> c0_n0_w7, 
            w8=> c0_n0_w8, 
            w9=> c0_n0_w9, 
            w10=> c0_n0_w10, 
            w11=> c0_n0_w11, 
            w12=> c0_n0_w12, 
            w13=> c0_n0_w13, 
            w14=> c0_n0_w14, 
            w15=> c0_n0_w15, 
            w16=> c0_n0_w16, 
            w17=> c0_n0_w17, 
            w18=> c0_n0_w18, 
            w19=> c0_n0_w19, 
            w20=> c0_n0_w20, 
            w21=> c0_n0_w21, 
            w22=> c0_n0_w22, 
            w23=> c0_n0_w23, 
            w24=> c0_n0_w24, 
            w25=> c0_n0_w25, 
            w26=> c0_n0_w26, 
            w27=> c0_n0_w27, 
            w28=> c0_n0_w28, 
            w29=> c0_n0_w29, 
            w30=> c0_n0_w30, 
            w31=> c0_n0_w31, 
            w32=> c0_n0_w32, 
            w33=> c0_n0_w33, 
            w34=> c0_n0_w34, 
            w35=> c0_n0_w35, 
            w36=> c0_n0_w36, 
            w37=> c0_n0_w37, 
            w38=> c0_n0_w38, 
            w39=> c0_n0_w39, 
            w40=> c0_n0_w40, 
            w41=> c0_n0_w41, 
            w42=> c0_n0_w42, 
            w43=> c0_n0_w43, 
            w44=> c0_n0_w44, 
            w45=> c0_n0_w45, 
            w46=> c0_n0_w46, 
            w47=> c0_n0_w47, 
            w48=> c0_n0_w48, 
            w49=> c0_n0_w49, 
            w50=> c0_n0_w50, 
            w51=> c0_n0_w51, 
            w52=> c0_n0_w52, 
            w53=> c0_n0_w53, 
            w54=> c0_n0_w54, 
            w55=> c0_n0_w55, 
            w56=> c0_n0_w56, 
            w57=> c0_n0_w57, 
            w58=> c0_n0_w58, 
            w59=> c0_n0_w59, 
            w60=> c0_n0_w60, 
            w61=> c0_n0_w61, 
            w62=> c0_n0_w62, 
            w63=> c0_n0_w63, 
            w64=> c0_n0_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n1_w1, 
            w2=> c0_n1_w2, 
            w3=> c0_n1_w3, 
            w4=> c0_n1_w4, 
            w5=> c0_n1_w5, 
            w6=> c0_n1_w6, 
            w7=> c0_n1_w7, 
            w8=> c0_n1_w8, 
            w9=> c0_n1_w9, 
            w10=> c0_n1_w10, 
            w11=> c0_n1_w11, 
            w12=> c0_n1_w12, 
            w13=> c0_n1_w13, 
            w14=> c0_n1_w14, 
            w15=> c0_n1_w15, 
            w16=> c0_n1_w16, 
            w17=> c0_n1_w17, 
            w18=> c0_n1_w18, 
            w19=> c0_n1_w19, 
            w20=> c0_n1_w20, 
            w21=> c0_n1_w21, 
            w22=> c0_n1_w22, 
            w23=> c0_n1_w23, 
            w24=> c0_n1_w24, 
            w25=> c0_n1_w25, 
            w26=> c0_n1_w26, 
            w27=> c0_n1_w27, 
            w28=> c0_n1_w28, 
            w29=> c0_n1_w29, 
            w30=> c0_n1_w30, 
            w31=> c0_n1_w31, 
            w32=> c0_n1_w32, 
            w33=> c0_n1_w33, 
            w34=> c0_n1_w34, 
            w35=> c0_n1_w35, 
            w36=> c0_n1_w36, 
            w37=> c0_n1_w37, 
            w38=> c0_n1_w38, 
            w39=> c0_n1_w39, 
            w40=> c0_n1_w40, 
            w41=> c0_n1_w41, 
            w42=> c0_n1_w42, 
            w43=> c0_n1_w43, 
            w44=> c0_n1_w44, 
            w45=> c0_n1_w45, 
            w46=> c0_n1_w46, 
            w47=> c0_n1_w47, 
            w48=> c0_n1_w48, 
            w49=> c0_n1_w49, 
            w50=> c0_n1_w50, 
            w51=> c0_n1_w51, 
            w52=> c0_n1_w52, 
            w53=> c0_n1_w53, 
            w54=> c0_n1_w54, 
            w55=> c0_n1_w55, 
            w56=> c0_n1_w56, 
            w57=> c0_n1_w57, 
            w58=> c0_n1_w58, 
            w59=> c0_n1_w59, 
            w60=> c0_n1_w60, 
            w61=> c0_n1_w61, 
            w62=> c0_n1_w62, 
            w63=> c0_n1_w63, 
            w64=> c0_n1_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n2_w1, 
            w2=> c0_n2_w2, 
            w3=> c0_n2_w3, 
            w4=> c0_n2_w4, 
            w5=> c0_n2_w5, 
            w6=> c0_n2_w6, 
            w7=> c0_n2_w7, 
            w8=> c0_n2_w8, 
            w9=> c0_n2_w9, 
            w10=> c0_n2_w10, 
            w11=> c0_n2_w11, 
            w12=> c0_n2_w12, 
            w13=> c0_n2_w13, 
            w14=> c0_n2_w14, 
            w15=> c0_n2_w15, 
            w16=> c0_n2_w16, 
            w17=> c0_n2_w17, 
            w18=> c0_n2_w18, 
            w19=> c0_n2_w19, 
            w20=> c0_n2_w20, 
            w21=> c0_n2_w21, 
            w22=> c0_n2_w22, 
            w23=> c0_n2_w23, 
            w24=> c0_n2_w24, 
            w25=> c0_n2_w25, 
            w26=> c0_n2_w26, 
            w27=> c0_n2_w27, 
            w28=> c0_n2_w28, 
            w29=> c0_n2_w29, 
            w30=> c0_n2_w30, 
            w31=> c0_n2_w31, 
            w32=> c0_n2_w32, 
            w33=> c0_n2_w33, 
            w34=> c0_n2_w34, 
            w35=> c0_n2_w35, 
            w36=> c0_n2_w36, 
            w37=> c0_n2_w37, 
            w38=> c0_n2_w38, 
            w39=> c0_n2_w39, 
            w40=> c0_n2_w40, 
            w41=> c0_n2_w41, 
            w42=> c0_n2_w42, 
            w43=> c0_n2_w43, 
            w44=> c0_n2_w44, 
            w45=> c0_n2_w45, 
            w46=> c0_n2_w46, 
            w47=> c0_n2_w47, 
            w48=> c0_n2_w48, 
            w49=> c0_n2_w49, 
            w50=> c0_n2_w50, 
            w51=> c0_n2_w51, 
            w52=> c0_n2_w52, 
            w53=> c0_n2_w53, 
            w54=> c0_n2_w54, 
            w55=> c0_n2_w55, 
            w56=> c0_n2_w56, 
            w57=> c0_n2_w57, 
            w58=> c0_n2_w58, 
            w59=> c0_n2_w59, 
            w60=> c0_n2_w60, 
            w61=> c0_n2_w61, 
            w62=> c0_n2_w62, 
            w63=> c0_n2_w63, 
            w64=> c0_n2_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n3_w1, 
            w2=> c0_n3_w2, 
            w3=> c0_n3_w3, 
            w4=> c0_n3_w4, 
            w5=> c0_n3_w5, 
            w6=> c0_n3_w6, 
            w7=> c0_n3_w7, 
            w8=> c0_n3_w8, 
            w9=> c0_n3_w9, 
            w10=> c0_n3_w10, 
            w11=> c0_n3_w11, 
            w12=> c0_n3_w12, 
            w13=> c0_n3_w13, 
            w14=> c0_n3_w14, 
            w15=> c0_n3_w15, 
            w16=> c0_n3_w16, 
            w17=> c0_n3_w17, 
            w18=> c0_n3_w18, 
            w19=> c0_n3_w19, 
            w20=> c0_n3_w20, 
            w21=> c0_n3_w21, 
            w22=> c0_n3_w22, 
            w23=> c0_n3_w23, 
            w24=> c0_n3_w24, 
            w25=> c0_n3_w25, 
            w26=> c0_n3_w26, 
            w27=> c0_n3_w27, 
            w28=> c0_n3_w28, 
            w29=> c0_n3_w29, 
            w30=> c0_n3_w30, 
            w31=> c0_n3_w31, 
            w32=> c0_n3_w32, 
            w33=> c0_n3_w33, 
            w34=> c0_n3_w34, 
            w35=> c0_n3_w35, 
            w36=> c0_n3_w36, 
            w37=> c0_n3_w37, 
            w38=> c0_n3_w38, 
            w39=> c0_n3_w39, 
            w40=> c0_n3_w40, 
            w41=> c0_n3_w41, 
            w42=> c0_n3_w42, 
            w43=> c0_n3_w43, 
            w44=> c0_n3_w44, 
            w45=> c0_n3_w45, 
            w46=> c0_n3_w46, 
            w47=> c0_n3_w47, 
            w48=> c0_n3_w48, 
            w49=> c0_n3_w49, 
            w50=> c0_n3_w50, 
            w51=> c0_n3_w51, 
            w52=> c0_n3_w52, 
            w53=> c0_n3_w53, 
            w54=> c0_n3_w54, 
            w55=> c0_n3_w55, 
            w56=> c0_n3_w56, 
            w57=> c0_n3_w57, 
            w58=> c0_n3_w58, 
            w59=> c0_n3_w59, 
            w60=> c0_n3_w60, 
            w61=> c0_n3_w61, 
            w62=> c0_n3_w62, 
            w63=> c0_n3_w63, 
            w64=> c0_n3_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n4_w1, 
            w2=> c0_n4_w2, 
            w3=> c0_n4_w3, 
            w4=> c0_n4_w4, 
            w5=> c0_n4_w5, 
            w6=> c0_n4_w6, 
            w7=> c0_n4_w7, 
            w8=> c0_n4_w8, 
            w9=> c0_n4_w9, 
            w10=> c0_n4_w10, 
            w11=> c0_n4_w11, 
            w12=> c0_n4_w12, 
            w13=> c0_n4_w13, 
            w14=> c0_n4_w14, 
            w15=> c0_n4_w15, 
            w16=> c0_n4_w16, 
            w17=> c0_n4_w17, 
            w18=> c0_n4_w18, 
            w19=> c0_n4_w19, 
            w20=> c0_n4_w20, 
            w21=> c0_n4_w21, 
            w22=> c0_n4_w22, 
            w23=> c0_n4_w23, 
            w24=> c0_n4_w24, 
            w25=> c0_n4_w25, 
            w26=> c0_n4_w26, 
            w27=> c0_n4_w27, 
            w28=> c0_n4_w28, 
            w29=> c0_n4_w29, 
            w30=> c0_n4_w30, 
            w31=> c0_n4_w31, 
            w32=> c0_n4_w32, 
            w33=> c0_n4_w33, 
            w34=> c0_n4_w34, 
            w35=> c0_n4_w35, 
            w36=> c0_n4_w36, 
            w37=> c0_n4_w37, 
            w38=> c0_n4_w38, 
            w39=> c0_n4_w39, 
            w40=> c0_n4_w40, 
            w41=> c0_n4_w41, 
            w42=> c0_n4_w42, 
            w43=> c0_n4_w43, 
            w44=> c0_n4_w44, 
            w45=> c0_n4_w45, 
            w46=> c0_n4_w46, 
            w47=> c0_n4_w47, 
            w48=> c0_n4_w48, 
            w49=> c0_n4_w49, 
            w50=> c0_n4_w50, 
            w51=> c0_n4_w51, 
            w52=> c0_n4_w52, 
            w53=> c0_n4_w53, 
            w54=> c0_n4_w54, 
            w55=> c0_n4_w55, 
            w56=> c0_n4_w56, 
            w57=> c0_n4_w57, 
            w58=> c0_n4_w58, 
            w59=> c0_n4_w59, 
            w60=> c0_n4_w60, 
            w61=> c0_n4_w61, 
            w62=> c0_n4_w62, 
            w63=> c0_n4_w63, 
            w64=> c0_n4_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n5_w1, 
            w2=> c0_n5_w2, 
            w3=> c0_n5_w3, 
            w4=> c0_n5_w4, 
            w5=> c0_n5_w5, 
            w6=> c0_n5_w6, 
            w7=> c0_n5_w7, 
            w8=> c0_n5_w8, 
            w9=> c0_n5_w9, 
            w10=> c0_n5_w10, 
            w11=> c0_n5_w11, 
            w12=> c0_n5_w12, 
            w13=> c0_n5_w13, 
            w14=> c0_n5_w14, 
            w15=> c0_n5_w15, 
            w16=> c0_n5_w16, 
            w17=> c0_n5_w17, 
            w18=> c0_n5_w18, 
            w19=> c0_n5_w19, 
            w20=> c0_n5_w20, 
            w21=> c0_n5_w21, 
            w22=> c0_n5_w22, 
            w23=> c0_n5_w23, 
            w24=> c0_n5_w24, 
            w25=> c0_n5_w25, 
            w26=> c0_n5_w26, 
            w27=> c0_n5_w27, 
            w28=> c0_n5_w28, 
            w29=> c0_n5_w29, 
            w30=> c0_n5_w30, 
            w31=> c0_n5_w31, 
            w32=> c0_n5_w32, 
            w33=> c0_n5_w33, 
            w34=> c0_n5_w34, 
            w35=> c0_n5_w35, 
            w36=> c0_n5_w36, 
            w37=> c0_n5_w37, 
            w38=> c0_n5_w38, 
            w39=> c0_n5_w39, 
            w40=> c0_n5_w40, 
            w41=> c0_n5_w41, 
            w42=> c0_n5_w42, 
            w43=> c0_n5_w43, 
            w44=> c0_n5_w44, 
            w45=> c0_n5_w45, 
            w46=> c0_n5_w46, 
            w47=> c0_n5_w47, 
            w48=> c0_n5_w48, 
            w49=> c0_n5_w49, 
            w50=> c0_n5_w50, 
            w51=> c0_n5_w51, 
            w52=> c0_n5_w52, 
            w53=> c0_n5_w53, 
            w54=> c0_n5_w54, 
            w55=> c0_n5_w55, 
            w56=> c0_n5_w56, 
            w57=> c0_n5_w57, 
            w58=> c0_n5_w58, 
            w59=> c0_n5_w59, 
            w60=> c0_n5_w60, 
            w61=> c0_n5_w61, 
            w62=> c0_n5_w62, 
            w63=> c0_n5_w63, 
            w64=> c0_n5_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n6_w1, 
            w2=> c0_n6_w2, 
            w3=> c0_n6_w3, 
            w4=> c0_n6_w4, 
            w5=> c0_n6_w5, 
            w6=> c0_n6_w6, 
            w7=> c0_n6_w7, 
            w8=> c0_n6_w8, 
            w9=> c0_n6_w9, 
            w10=> c0_n6_w10, 
            w11=> c0_n6_w11, 
            w12=> c0_n6_w12, 
            w13=> c0_n6_w13, 
            w14=> c0_n6_w14, 
            w15=> c0_n6_w15, 
            w16=> c0_n6_w16, 
            w17=> c0_n6_w17, 
            w18=> c0_n6_w18, 
            w19=> c0_n6_w19, 
            w20=> c0_n6_w20, 
            w21=> c0_n6_w21, 
            w22=> c0_n6_w22, 
            w23=> c0_n6_w23, 
            w24=> c0_n6_w24, 
            w25=> c0_n6_w25, 
            w26=> c0_n6_w26, 
            w27=> c0_n6_w27, 
            w28=> c0_n6_w28, 
            w29=> c0_n6_w29, 
            w30=> c0_n6_w30, 
            w31=> c0_n6_w31, 
            w32=> c0_n6_w32, 
            w33=> c0_n6_w33, 
            w34=> c0_n6_w34, 
            w35=> c0_n6_w35, 
            w36=> c0_n6_w36, 
            w37=> c0_n6_w37, 
            w38=> c0_n6_w38, 
            w39=> c0_n6_w39, 
            w40=> c0_n6_w40, 
            w41=> c0_n6_w41, 
            w42=> c0_n6_w42, 
            w43=> c0_n6_w43, 
            w44=> c0_n6_w44, 
            w45=> c0_n6_w45, 
            w46=> c0_n6_w46, 
            w47=> c0_n6_w47, 
            w48=> c0_n6_w48, 
            w49=> c0_n6_w49, 
            w50=> c0_n6_w50, 
            w51=> c0_n6_w51, 
            w52=> c0_n6_w52, 
            w53=> c0_n6_w53, 
            w54=> c0_n6_w54, 
            w55=> c0_n6_w55, 
            w56=> c0_n6_w56, 
            w57=> c0_n6_w57, 
            w58=> c0_n6_w58, 
            w59=> c0_n6_w59, 
            w60=> c0_n6_w60, 
            w61=> c0_n6_w61, 
            w62=> c0_n6_w62, 
            w63=> c0_n6_w63, 
            w64=> c0_n6_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n7_w1, 
            w2=> c0_n7_w2, 
            w3=> c0_n7_w3, 
            w4=> c0_n7_w4, 
            w5=> c0_n7_w5, 
            w6=> c0_n7_w6, 
            w7=> c0_n7_w7, 
            w8=> c0_n7_w8, 
            w9=> c0_n7_w9, 
            w10=> c0_n7_w10, 
            w11=> c0_n7_w11, 
            w12=> c0_n7_w12, 
            w13=> c0_n7_w13, 
            w14=> c0_n7_w14, 
            w15=> c0_n7_w15, 
            w16=> c0_n7_w16, 
            w17=> c0_n7_w17, 
            w18=> c0_n7_w18, 
            w19=> c0_n7_w19, 
            w20=> c0_n7_w20, 
            w21=> c0_n7_w21, 
            w22=> c0_n7_w22, 
            w23=> c0_n7_w23, 
            w24=> c0_n7_w24, 
            w25=> c0_n7_w25, 
            w26=> c0_n7_w26, 
            w27=> c0_n7_w27, 
            w28=> c0_n7_w28, 
            w29=> c0_n7_w29, 
            w30=> c0_n7_w30, 
            w31=> c0_n7_w31, 
            w32=> c0_n7_w32, 
            w33=> c0_n7_w33, 
            w34=> c0_n7_w34, 
            w35=> c0_n7_w35, 
            w36=> c0_n7_w36, 
            w37=> c0_n7_w37, 
            w38=> c0_n7_w38, 
            w39=> c0_n7_w39, 
            w40=> c0_n7_w40, 
            w41=> c0_n7_w41, 
            w42=> c0_n7_w42, 
            w43=> c0_n7_w43, 
            w44=> c0_n7_w44, 
            w45=> c0_n7_w45, 
            w46=> c0_n7_w46, 
            w47=> c0_n7_w47, 
            w48=> c0_n7_w48, 
            w49=> c0_n7_w49, 
            w50=> c0_n7_w50, 
            w51=> c0_n7_w51, 
            w52=> c0_n7_w52, 
            w53=> c0_n7_w53, 
            w54=> c0_n7_w54, 
            w55=> c0_n7_w55, 
            w56=> c0_n7_w56, 
            w57=> c0_n7_w57, 
            w58=> c0_n7_w58, 
            w59=> c0_n7_w59, 
            w60=> c0_n7_w60, 
            w61=> c0_n7_w61, 
            w62=> c0_n7_w62, 
            w63=> c0_n7_w63, 
            w64=> c0_n7_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n8_w1, 
            w2=> c0_n8_w2, 
            w3=> c0_n8_w3, 
            w4=> c0_n8_w4, 
            w5=> c0_n8_w5, 
            w6=> c0_n8_w6, 
            w7=> c0_n8_w7, 
            w8=> c0_n8_w8, 
            w9=> c0_n8_w9, 
            w10=> c0_n8_w10, 
            w11=> c0_n8_w11, 
            w12=> c0_n8_w12, 
            w13=> c0_n8_w13, 
            w14=> c0_n8_w14, 
            w15=> c0_n8_w15, 
            w16=> c0_n8_w16, 
            w17=> c0_n8_w17, 
            w18=> c0_n8_w18, 
            w19=> c0_n8_w19, 
            w20=> c0_n8_w20, 
            w21=> c0_n8_w21, 
            w22=> c0_n8_w22, 
            w23=> c0_n8_w23, 
            w24=> c0_n8_w24, 
            w25=> c0_n8_w25, 
            w26=> c0_n8_w26, 
            w27=> c0_n8_w27, 
            w28=> c0_n8_w28, 
            w29=> c0_n8_w29, 
            w30=> c0_n8_w30, 
            w31=> c0_n8_w31, 
            w32=> c0_n8_w32, 
            w33=> c0_n8_w33, 
            w34=> c0_n8_w34, 
            w35=> c0_n8_w35, 
            w36=> c0_n8_w36, 
            w37=> c0_n8_w37, 
            w38=> c0_n8_w38, 
            w39=> c0_n8_w39, 
            w40=> c0_n8_w40, 
            w41=> c0_n8_w41, 
            w42=> c0_n8_w42, 
            w43=> c0_n8_w43, 
            w44=> c0_n8_w44, 
            w45=> c0_n8_w45, 
            w46=> c0_n8_w46, 
            w47=> c0_n8_w47, 
            w48=> c0_n8_w48, 
            w49=> c0_n8_w49, 
            w50=> c0_n8_w50, 
            w51=> c0_n8_w51, 
            w52=> c0_n8_w52, 
            w53=> c0_n8_w53, 
            w54=> c0_n8_w54, 
            w55=> c0_n8_w55, 
            w56=> c0_n8_w56, 
            w57=> c0_n8_w57, 
            w58=> c0_n8_w58, 
            w59=> c0_n8_w59, 
            w60=> c0_n8_w60, 
            w61=> c0_n8_w61, 
            w62=> c0_n8_w62, 
            w63=> c0_n8_w63, 
            w64=> c0_n8_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n9_w1, 
            w2=> c0_n9_w2, 
            w3=> c0_n9_w3, 
            w4=> c0_n9_w4, 
            w5=> c0_n9_w5, 
            w6=> c0_n9_w6, 
            w7=> c0_n9_w7, 
            w8=> c0_n9_w8, 
            w9=> c0_n9_w9, 
            w10=> c0_n9_w10, 
            w11=> c0_n9_w11, 
            w12=> c0_n9_w12, 
            w13=> c0_n9_w13, 
            w14=> c0_n9_w14, 
            w15=> c0_n9_w15, 
            w16=> c0_n9_w16, 
            w17=> c0_n9_w17, 
            w18=> c0_n9_w18, 
            w19=> c0_n9_w19, 
            w20=> c0_n9_w20, 
            w21=> c0_n9_w21, 
            w22=> c0_n9_w22, 
            w23=> c0_n9_w23, 
            w24=> c0_n9_w24, 
            w25=> c0_n9_w25, 
            w26=> c0_n9_w26, 
            w27=> c0_n9_w27, 
            w28=> c0_n9_w28, 
            w29=> c0_n9_w29, 
            w30=> c0_n9_w30, 
            w31=> c0_n9_w31, 
            w32=> c0_n9_w32, 
            w33=> c0_n9_w33, 
            w34=> c0_n9_w34, 
            w35=> c0_n9_w35, 
            w36=> c0_n9_w36, 
            w37=> c0_n9_w37, 
            w38=> c0_n9_w38, 
            w39=> c0_n9_w39, 
            w40=> c0_n9_w40, 
            w41=> c0_n9_w41, 
            w42=> c0_n9_w42, 
            w43=> c0_n9_w43, 
            w44=> c0_n9_w44, 
            w45=> c0_n9_w45, 
            w46=> c0_n9_w46, 
            w47=> c0_n9_w47, 
            w48=> c0_n9_w48, 
            w49=> c0_n9_w49, 
            w50=> c0_n9_w50, 
            w51=> c0_n9_w51, 
            w52=> c0_n9_w52, 
            w53=> c0_n9_w53, 
            w54=> c0_n9_w54, 
            w55=> c0_n9_w55, 
            w56=> c0_n9_w56, 
            w57=> c0_n9_w57, 
            w58=> c0_n9_w58, 
            w59=> c0_n9_w59, 
            w60=> c0_n9_w60, 
            w61=> c0_n9_w61, 
            w62=> c0_n9_w62, 
            w63=> c0_n9_w63, 
            w64=> c0_n9_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n9_y
   );           
            
neuron_inst_10: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n10_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n10_w1, 
            w2=> c0_n10_w2, 
            w3=> c0_n10_w3, 
            w4=> c0_n10_w4, 
            w5=> c0_n10_w5, 
            w6=> c0_n10_w6, 
            w7=> c0_n10_w7, 
            w8=> c0_n10_w8, 
            w9=> c0_n10_w9, 
            w10=> c0_n10_w10, 
            w11=> c0_n10_w11, 
            w12=> c0_n10_w12, 
            w13=> c0_n10_w13, 
            w14=> c0_n10_w14, 
            w15=> c0_n10_w15, 
            w16=> c0_n10_w16, 
            w17=> c0_n10_w17, 
            w18=> c0_n10_w18, 
            w19=> c0_n10_w19, 
            w20=> c0_n10_w20, 
            w21=> c0_n10_w21, 
            w22=> c0_n10_w22, 
            w23=> c0_n10_w23, 
            w24=> c0_n10_w24, 
            w25=> c0_n10_w25, 
            w26=> c0_n10_w26, 
            w27=> c0_n10_w27, 
            w28=> c0_n10_w28, 
            w29=> c0_n10_w29, 
            w30=> c0_n10_w30, 
            w31=> c0_n10_w31, 
            w32=> c0_n10_w32, 
            w33=> c0_n10_w33, 
            w34=> c0_n10_w34, 
            w35=> c0_n10_w35, 
            w36=> c0_n10_w36, 
            w37=> c0_n10_w37, 
            w38=> c0_n10_w38, 
            w39=> c0_n10_w39, 
            w40=> c0_n10_w40, 
            w41=> c0_n10_w41, 
            w42=> c0_n10_w42, 
            w43=> c0_n10_w43, 
            w44=> c0_n10_w44, 
            w45=> c0_n10_w45, 
            w46=> c0_n10_w46, 
            w47=> c0_n10_w47, 
            w48=> c0_n10_w48, 
            w49=> c0_n10_w49, 
            w50=> c0_n10_w50, 
            w51=> c0_n10_w51, 
            w52=> c0_n10_w52, 
            w53=> c0_n10_w53, 
            w54=> c0_n10_w54, 
            w55=> c0_n10_w55, 
            w56=> c0_n10_w56, 
            w57=> c0_n10_w57, 
            w58=> c0_n10_w58, 
            w59=> c0_n10_w59, 
            w60=> c0_n10_w60, 
            w61=> c0_n10_w61, 
            w62=> c0_n10_w62, 
            w63=> c0_n10_w63, 
            w64=> c0_n10_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n10_y
   );           
            
neuron_inst_11: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n11_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n11_w1, 
            w2=> c0_n11_w2, 
            w3=> c0_n11_w3, 
            w4=> c0_n11_w4, 
            w5=> c0_n11_w5, 
            w6=> c0_n11_w6, 
            w7=> c0_n11_w7, 
            w8=> c0_n11_w8, 
            w9=> c0_n11_w9, 
            w10=> c0_n11_w10, 
            w11=> c0_n11_w11, 
            w12=> c0_n11_w12, 
            w13=> c0_n11_w13, 
            w14=> c0_n11_w14, 
            w15=> c0_n11_w15, 
            w16=> c0_n11_w16, 
            w17=> c0_n11_w17, 
            w18=> c0_n11_w18, 
            w19=> c0_n11_w19, 
            w20=> c0_n11_w20, 
            w21=> c0_n11_w21, 
            w22=> c0_n11_w22, 
            w23=> c0_n11_w23, 
            w24=> c0_n11_w24, 
            w25=> c0_n11_w25, 
            w26=> c0_n11_w26, 
            w27=> c0_n11_w27, 
            w28=> c0_n11_w28, 
            w29=> c0_n11_w29, 
            w30=> c0_n11_w30, 
            w31=> c0_n11_w31, 
            w32=> c0_n11_w32, 
            w33=> c0_n11_w33, 
            w34=> c0_n11_w34, 
            w35=> c0_n11_w35, 
            w36=> c0_n11_w36, 
            w37=> c0_n11_w37, 
            w38=> c0_n11_w38, 
            w39=> c0_n11_w39, 
            w40=> c0_n11_w40, 
            w41=> c0_n11_w41, 
            w42=> c0_n11_w42, 
            w43=> c0_n11_w43, 
            w44=> c0_n11_w44, 
            w45=> c0_n11_w45, 
            w46=> c0_n11_w46, 
            w47=> c0_n11_w47, 
            w48=> c0_n11_w48, 
            w49=> c0_n11_w49, 
            w50=> c0_n11_w50, 
            w51=> c0_n11_w51, 
            w52=> c0_n11_w52, 
            w53=> c0_n11_w53, 
            w54=> c0_n11_w54, 
            w55=> c0_n11_w55, 
            w56=> c0_n11_w56, 
            w57=> c0_n11_w57, 
            w58=> c0_n11_w58, 
            w59=> c0_n11_w59, 
            w60=> c0_n11_w60, 
            w61=> c0_n11_w61, 
            w62=> c0_n11_w62, 
            w63=> c0_n11_w63, 
            w64=> c0_n11_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n11_y
   );           
            
neuron_inst_12: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n12_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n12_w1, 
            w2=> c0_n12_w2, 
            w3=> c0_n12_w3, 
            w4=> c0_n12_w4, 
            w5=> c0_n12_w5, 
            w6=> c0_n12_w6, 
            w7=> c0_n12_w7, 
            w8=> c0_n12_w8, 
            w9=> c0_n12_w9, 
            w10=> c0_n12_w10, 
            w11=> c0_n12_w11, 
            w12=> c0_n12_w12, 
            w13=> c0_n12_w13, 
            w14=> c0_n12_w14, 
            w15=> c0_n12_w15, 
            w16=> c0_n12_w16, 
            w17=> c0_n12_w17, 
            w18=> c0_n12_w18, 
            w19=> c0_n12_w19, 
            w20=> c0_n12_w20, 
            w21=> c0_n12_w21, 
            w22=> c0_n12_w22, 
            w23=> c0_n12_w23, 
            w24=> c0_n12_w24, 
            w25=> c0_n12_w25, 
            w26=> c0_n12_w26, 
            w27=> c0_n12_w27, 
            w28=> c0_n12_w28, 
            w29=> c0_n12_w29, 
            w30=> c0_n12_w30, 
            w31=> c0_n12_w31, 
            w32=> c0_n12_w32, 
            w33=> c0_n12_w33, 
            w34=> c0_n12_w34, 
            w35=> c0_n12_w35, 
            w36=> c0_n12_w36, 
            w37=> c0_n12_w37, 
            w38=> c0_n12_w38, 
            w39=> c0_n12_w39, 
            w40=> c0_n12_w40, 
            w41=> c0_n12_w41, 
            w42=> c0_n12_w42, 
            w43=> c0_n12_w43, 
            w44=> c0_n12_w44, 
            w45=> c0_n12_w45, 
            w46=> c0_n12_w46, 
            w47=> c0_n12_w47, 
            w48=> c0_n12_w48, 
            w49=> c0_n12_w49, 
            w50=> c0_n12_w50, 
            w51=> c0_n12_w51, 
            w52=> c0_n12_w52, 
            w53=> c0_n12_w53, 
            w54=> c0_n12_w54, 
            w55=> c0_n12_w55, 
            w56=> c0_n12_w56, 
            w57=> c0_n12_w57, 
            w58=> c0_n12_w58, 
            w59=> c0_n12_w59, 
            w60=> c0_n12_w60, 
            w61=> c0_n12_w61, 
            w62=> c0_n12_w62, 
            w63=> c0_n12_w63, 
            w64=> c0_n12_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n12_y
   );           
            
neuron_inst_13: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n13_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n13_w1, 
            w2=> c0_n13_w2, 
            w3=> c0_n13_w3, 
            w4=> c0_n13_w4, 
            w5=> c0_n13_w5, 
            w6=> c0_n13_w6, 
            w7=> c0_n13_w7, 
            w8=> c0_n13_w8, 
            w9=> c0_n13_w9, 
            w10=> c0_n13_w10, 
            w11=> c0_n13_w11, 
            w12=> c0_n13_w12, 
            w13=> c0_n13_w13, 
            w14=> c0_n13_w14, 
            w15=> c0_n13_w15, 
            w16=> c0_n13_w16, 
            w17=> c0_n13_w17, 
            w18=> c0_n13_w18, 
            w19=> c0_n13_w19, 
            w20=> c0_n13_w20, 
            w21=> c0_n13_w21, 
            w22=> c0_n13_w22, 
            w23=> c0_n13_w23, 
            w24=> c0_n13_w24, 
            w25=> c0_n13_w25, 
            w26=> c0_n13_w26, 
            w27=> c0_n13_w27, 
            w28=> c0_n13_w28, 
            w29=> c0_n13_w29, 
            w30=> c0_n13_w30, 
            w31=> c0_n13_w31, 
            w32=> c0_n13_w32, 
            w33=> c0_n13_w33, 
            w34=> c0_n13_w34, 
            w35=> c0_n13_w35, 
            w36=> c0_n13_w36, 
            w37=> c0_n13_w37, 
            w38=> c0_n13_w38, 
            w39=> c0_n13_w39, 
            w40=> c0_n13_w40, 
            w41=> c0_n13_w41, 
            w42=> c0_n13_w42, 
            w43=> c0_n13_w43, 
            w44=> c0_n13_w44, 
            w45=> c0_n13_w45, 
            w46=> c0_n13_w46, 
            w47=> c0_n13_w47, 
            w48=> c0_n13_w48, 
            w49=> c0_n13_w49, 
            w50=> c0_n13_w50, 
            w51=> c0_n13_w51, 
            w52=> c0_n13_w52, 
            w53=> c0_n13_w53, 
            w54=> c0_n13_w54, 
            w55=> c0_n13_w55, 
            w56=> c0_n13_w56, 
            w57=> c0_n13_w57, 
            w58=> c0_n13_w58, 
            w59=> c0_n13_w59, 
            w60=> c0_n13_w60, 
            w61=> c0_n13_w61, 
            w62=> c0_n13_w62, 
            w63=> c0_n13_w63, 
            w64=> c0_n13_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n13_y
   );           
            
neuron_inst_14: ENTITY work.neuron_comb_ReLU_64n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n14_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            w1=> c0_n14_w1, 
            w2=> c0_n14_w2, 
            w3=> c0_n14_w3, 
            w4=> c0_n14_w4, 
            w5=> c0_n14_w5, 
            w6=> c0_n14_w6, 
            w7=> c0_n14_w7, 
            w8=> c0_n14_w8, 
            w9=> c0_n14_w9, 
            w10=> c0_n14_w10, 
            w11=> c0_n14_w11, 
            w12=> c0_n14_w12, 
            w13=> c0_n14_w13, 
            w14=> c0_n14_w14, 
            w15=> c0_n14_w15, 
            w16=> c0_n14_w16, 
            w17=> c0_n14_w17, 
            w18=> c0_n14_w18, 
            w19=> c0_n14_w19, 
            w20=> c0_n14_w20, 
            w21=> c0_n14_w21, 
            w22=> c0_n14_w22, 
            w23=> c0_n14_w23, 
            w24=> c0_n14_w24, 
            w25=> c0_n14_w25, 
            w26=> c0_n14_w26, 
            w27=> c0_n14_w27, 
            w28=> c0_n14_w28, 
            w29=> c0_n14_w29, 
            w30=> c0_n14_w30, 
            w31=> c0_n14_w31, 
            w32=> c0_n14_w32, 
            w33=> c0_n14_w33, 
            w34=> c0_n14_w34, 
            w35=> c0_n14_w35, 
            w36=> c0_n14_w36, 
            w37=> c0_n14_w37, 
            w38=> c0_n14_w38, 
            w39=> c0_n14_w39, 
            w40=> c0_n14_w40, 
            w41=> c0_n14_w41, 
            w42=> c0_n14_w42, 
            w43=> c0_n14_w43, 
            w44=> c0_n14_w44, 
            w45=> c0_n14_w45, 
            w46=> c0_n14_w46, 
            w47=> c0_n14_w47, 
            w48=> c0_n14_w48, 
            w49=> c0_n14_w49, 
            w50=> c0_n14_w50, 
            w51=> c0_n14_w51, 
            w52=> c0_n14_w52, 
            w53=> c0_n14_w53, 
            w54=> c0_n14_w54, 
            w55=> c0_n14_w55, 
            w56=> c0_n14_w56, 
            w57=> c0_n14_w57, 
            w58=> c0_n14_w58, 
            w59=> c0_n14_w59, 
            w60=> c0_n14_w60, 
            w61=> c0_n14_w61, 
            w62=> c0_n14_w62, 
            w63=> c0_n14_w63, 
            w64=> c0_n14_w64, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n14_y
   );           
             
END ARCHITECTURE;
