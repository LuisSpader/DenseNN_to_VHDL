
--https://stackoverflow.com/questions/17579716/implementing-rom-in-xilinx-vhdl
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.numeric_std.all;
----------------
ENTITY ROM_fx_10bitaddr_10width is
generic(addr_heigth : integer := 1024; -- store 1024 elements
				addr_bits  : integer := 10; -- required bits to store 1024 elements
				data_width : integer := 10  -- each element has 10-bits
				);
  PORT (
    address : IN STD_LOGIC_VECTOR(addr_bits - 1 DOWNTO 0);
    data_out : OUT STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0)
  );
END ENTITY;
------------------
architecture arch of ROM_fx_10bitaddr_10width is
	type memory is array ( 0 to addr_heigth-1 ) of std_logic_vector(data_width-1 downto 0 ) ;
	constant myrom : memory := (
--"int_f_x",--(address)  =integer_MAC|| f(x)               = int_f_x 
"1000000000",-- (0000000000) = 0.0       || 512.0              = 512.0
"1000000010",-- (0000000001) = 1.0       || 514.7999720869225  = 514.0
"1000000101",-- (0000000010) = 2.0       || 517.5997767033934  = 517.0
"1000001000",-- (0000000011) = 3.0       || 520.3992464190255  = 520.0
"1000001011",-- (0000000100) = 4.0       || 523.1982138835398  = 523.0
"1000001101",-- (0000000101) = 5.0       || 525.996511866768   = 525.0
"1000010000",-- (0000000110) = 6.0       || 528.7939732985955  = 528.0
"1000010011",-- (0000000111) = 7.0       || 531.5904313088217  = 531.0
"1000010110",-- (0000001000) = 8.0       || 534.38571926692    = 534.0
"1000011001",-- (0000001001) = 9.0       || 537.1796708216743  = 537.0
"1000011011",-- (0000001010) = 10.0      || 539.9721199406767  = 539.0
"1000011110",-- (0000001011) = 11.0      || 542.7629009496613  = 542.0
"1000100001",-- (0000001100) = 12.0      || 545.5518485716582  = 545.0
"1000100100",-- (0000001101) = 13.0      || 548.3387979659461  = 548.0
"1000100111",-- (0000001110) = 14.0      || 551.1235847667854  = 551.0
"1000101001",-- (0000001111) = 15.0      || 553.9060451219113  = 553.0
"1000101100",-- (0000010000) = 16.0      || 556.6860157307688  = 556.0
"1000101111",-- (0000010001) = 17.0      || 559.4633338824706  = 559.0
"1000110010",-- (0000010010) = 18.0      || 562.2378374934598  = 562.0
"1000110101",-- (0000010011) = 19.0      || 565.0093651448569  = 565.0
"1000110111",-- (0000010100) = 20.0      || 567.7777561194775  = 567.0
"1000111010",-- (0000010101) = 21.0      || 570.5428504384977  = 570.0
"1000111101",-- (0000010110) = 22.0      || 573.3044888977539  = 573.0
"1001000000",-- (0000010111) = 23.0      || 576.0625131036578  = 576.0
"1001000010",-- (0000011000) = 24.0      || 578.8167655087103  = 578.0
"1001000101",-- (0000011001) = 25.0      || 581.567089446598   = 581.0
"1001001000",-- (0000011010) = 26.0      || 584.3133291668554  = 584.0
"1001001011",-- (0000011011) = 27.0      || 587.055329869079   = 587.0
"1001001101",-- (0000011100) = 28.0      || 589.792937736675   = 589.0
"1001010000",-- (0000011101) = 29.0      || 592.5259999701284  = 592.0
"1001010011",-- (0000011110) = 30.0      || 595.2543648197768  = 595.0
"1001010101",-- (0000011111) = 31.0      || 597.9778816180766  = 597.0
"1001011000",-- (0000100000) = 32.0      || 600.696400811346   = 600.0
"1001011011",-- (0000100001) = 33.0      || 603.4097739909726  = 603.0
"1001011110",-- (0000100010) = 34.0      || 606.1178539240724  = 606.0
"1001100000",-- (0000100011) = 35.0      || 608.8204945835885  = 608.0
"1001100011",-- (0000100100) = 36.0      || 611.5175511778144  = 611.0
"1001100110",-- (0000100101) = 37.0      || 614.2088801793358  = 614.0
"1001101000",-- (0000100110) = 38.0      || 616.8943393533742  = 616.0
"1001101011",-- (0000100111) = 39.0      || 619.5737877855254  = 619.0
"1001101110",-- (0000101000) = 40.0      || 622.2470859088811  = 622.0
"1001110000",-- (0000101001) = 41.0      || 624.9140955305239  = 624.0
"1001110011",-- (0000101010) = 42.0      || 627.5746798573888  = 627.0
"1001110110",-- (0000101011) = 43.0      || 630.2287035214774  = 630.0
"1001111000",-- (0000101100) = 44.0      || 632.8760326044237  = 632.0
"1001111011",-- (0000101101) = 45.0      || 635.5165346613968  = 635.0
"1001111110",-- (0000101110) = 46.0      || 638.1500787443384  = 638.0
"1010000000",-- (0000101111) = 47.0      || 640.7765354245258  = 640.0
"1010000011",-- (0000110000) = 48.0      || 643.3957768144551  = 643.0
"1010000110",-- (0000110001) = 49.0      || 646.0076765890378  = 646.0
"1010001000",-- (0000110010) = 50.0      || 648.6121100061083  = 648.0
"1010001011",-- (0000110011) = 51.0      || 651.2089539262341  = 651.0
"1010001101",-- (0000110100) = 52.0      || 653.7980868318268  = 653.0
"1010010000",-- (0000110101) = 53.0      || 656.3793888455496  = 656.0
"1010010010",-- (0000110110) = 54.0      || 658.9527417480184  = 658.0
"1010010101",-- (0000110111) = 55.0      || 661.5180289947925  = 661.0
"1010011000",-- (0000111000) = 56.0      || 664.075135732655   = 664.0
"1010011010",-- (0000111001) = 57.0      || 666.6239488151787  = 666.0
"1010011101",-- (0000111010) = 58.0      || 669.1643568175771  = 669.0
"1010011111",-- (0000111011) = 59.0      || 671.6962500508422  = 671.0
"1010100010",-- (0000111100) = 60.0      || 674.2195205751634  = 674.0
"1010100100",-- (0000111101) = 61.0      || 676.7340622126334  = 676.0
"1010100111",-- (0000111110) = 62.0      || 679.2397705592377  = 679.0
"1010101001",-- (0000111111) = 63.0      || 681.7365429961313  = 681.0
"1010101100",-- (0001000000) = 64.0      || 684.2242787002021  = 684.0
"1010101110",-- (0001000001) = 65.0      || 686.7028786539244  = 686.0
"1010110001",-- (0001000010) = 66.0      || 689.1722456545049  = 689.0
"1010110011",-- (0001000011) = 67.0      || 691.6322843223231  = 691.0
"1010110110",-- (0001000100) = 68.0      || 694.0829011086701  = 694.0
"1010111000",-- (0001000101) = 69.0      || 696.5240043027885  = 696.0
"1010111010",-- (0001000110) = 70.0      || 698.9555040382198  = 698.0
"1010111101",-- (0001000111) = 71.0      || 701.3773122984612  = 701.0
"1010111111",-- (0001001000) = 72.0      || 703.7893429219371  = 703.0
"1011000010",-- (0001001001) = 73.0      || 706.1915116062916  = 706.0
"1011000100",-- (0001001010) = 74.0      || 708.5837359120085  = 708.0
"1011000110",-- (0001001011) = 75.0      || 710.9659352653605  = 710.0
"1011001001",-- (0001001100) = 76.0      || 713.3380309606988  = 713.0
"1011001011",-- (0001001101) = 77.0      || 715.6999461620873  = 715.0
"1011001110",-- (0001001110) = 78.0      || 718.0516059042876  = 718.0
"1011010000",-- (0001001111) = 79.0      || 720.392937093105   = 720.0
"1011010010",-- (0001010000) = 80.0      || 722.7238685050995  = 722.0
"1011010101",-- (0001010001) = 81.0      || 725.0443307866723  = 725.0
"1011010111",-- (0001010010) = 82.0      || 727.354256452535   = 727.0
"1011011001",-- (0001010011) = 83.0      || 729.6535798835699  = 729.0
"1011011011",-- (0001010100) = 84.0      || 731.9422373240906  = 731.0
"1011011110",-- (0001010101) = 85.0      || 734.2201668785095  = 734.0
"1011100000",-- (0001010110) = 86.0      || 736.4873085074267  = 736.0
"1011100010",-- (0001010111) = 87.0      || 738.7436040231428  = 738.0
"1011100100",-- (0001011000) = 88.0      || 740.9889970846107  = 740.0
"1011100111",-- (0001011001) = 89.0      || 743.223433191834   = 743.0
"1011101001",-- (0001011010) = 90.0      || 745.4468596797209  = 745.0
"1011101011",-- (0001011011) = 91.0      || 747.6592257114072  = 747.0
"1011101101",-- (0001011100) = 92.0      || 749.8604822710545  = 749.0
"1011110000",-- (0001011101) = 93.0      || 752.0505821561377  = 752.0
"1011110010",-- (0001011110) = 94.0      || 754.229479969231   = 754.0
"1011110100",-- (0001011111) = 95.0      || 756.3971321093014  = 756.0
"1011110110",-- (0001100000) = 96.0      || 758.5534967625256  = 758.0
"1011111000",-- (0001100001) = 97.0      || 760.6985338926354  = 760.0
"1011111010",-- (0001100010) = 98.0      || 762.8322052308068  = 762.0
"1011111100",-- (0001100011) = 99.0      || 764.9544742651028  = 764.0
"1011111111",-- (0001100100) = 100.0     || 767.0653062294809  = 767.0
"1100000001",-- (0001100101) = 101.0     || 769.1646680923774  = 769.0
"1100000011",-- (0001100110) = 102.0     || 771.252528544879   = 771.0
"1100000101",-- (0001100111) = 103.0     || 773.3288579884944  = 773.0
"1100000111",-- (0001101000) = 104.0     || 775.3936285225369  = 775.0
"1100001001",-- (0001101001) = 105.0     || 777.4468139311285  = 777.0
"1100001011",-- (0001101010) = 106.0     || 779.4883896698399  = 779.0
"1100001101",-- (0001101011) = 107.0     || 781.5183328519739  = 781.0
"1100001111",-- (0001101100) = 108.0     || 783.5366222345098  = 783.0
"1100010001",-- (0001101101) = 109.0     || 785.5432382037125  = 785.0
"1100010011",-- (0001101110) = 110.0     || 787.5381627604257  = 787.0
"1100010101",-- (0001101111) = 111.0     || 789.5213795050558  = 789.0
"1100010111",-- (0001110000) = 112.0     || 791.4928736222603  = 791.0
"1100011001",-- (0001110001) = 113.0     || 793.4526318653504  = 793.0
"1100011011",-- (0001110010) = 114.0     || 795.4006425404219  = 795.0
"1100011101",-- (0001110011) = 115.0     || 797.3368954902243  = 797.0
"1100011111",-- (0001110100) = 116.0     || 799.2613820777768  = 799.0
"1100100001",-- (0001110101) = 117.0     || 801.1740951697506  = 801.0
"1100100011",-- (0001110110) = 118.0     || 803.0750291196168  = 803.0
"1100100100",-- (0001110111) = 119.0     || 804.9641797505838  = 804.0
"1100100110",-- (0001111000) = 120.0     || 806.8415443383242  = 806.0
"1100101000",-- (0001111001) = 121.0     || 808.7071215935099  = 808.0
"1100101010",-- (0001111010) = 122.0     || 810.560911644163   = 810.0
"1100101100",-- (0001111011) = 123.0     || 812.4029160178314  = 812.0
"1100101110",-- (0001111100) = 124.0     || 814.2331376236062  = 814.0
"1100110000",-- (0001111101) = 125.0     || 816.0515807339825  = 816.0
"1100110001",-- (0001111110) = 126.0     || 817.8582509665817  = 817.0
"1100110011",-- (0001111111) = 127.0     || 819.6531552657422  = 819.0
"1100110101",-- (0010000000) = 128.0     || 821.4363018839877  = 821.0
"1100110111",-- (0010000001) = 129.0     || 823.207700363386   = 823.0
"1100111000",-- (0010000010) = 130.0     || 824.9673615168055  = 824.0
"1100111010",-- (0010000011) = 131.0     || 826.7152974090802  = 826.0
"1100111100",-- (0010000100) = 132.0     || 828.4515213380944  = 828.0
"1100111110",-- (0010000101) = 133.0     || 830.1760478157914  = 830.0
"1100111111",-- (0010000110) = 134.0     || 831.8888925491236  = 831.0
"1101000001",-- (0010000111) = 135.0     || 833.5900724209442  = 833.0
"1101000011",-- (0010001000) = 136.0     || 835.279605470856   = 835.0
"1101000100",-- (0010001001) = 137.0     || 836.9575108760243  = 836.0
"1101000110",-- (0010001010) = 138.0     || 838.623808931959   = 838.0
"1101001000",-- (0010001011) = 139.0     || 840.2785210332817  = 840.0
"1101001001",-- (0010001100) = 140.0     || 841.9216696544771  = 841.0
"1101001011",-- (0010001101) = 141.0     || 843.5532783306461  = 843.0
"1101001101",-- (0010001110) = 142.0     || 845.1733716382595  = 845.0
"1101001110",-- (0010001111) = 143.0     || 846.7819751759279  = 846.0
"1101010000",-- (0010010000) = 144.0     || 848.3791155451895  = 848.0
"1101010001",-- (0010010001) = 145.0     || 849.9648203313279  = 849.0
"1101010011",-- (0010010010) = 146.0     || 851.5391180842223  = 851.0
"1101010101",-- (0010010011) = 147.0     || 853.1020382992426  = 853.0
"1101010110",-- (0010010100) = 148.0     || 854.6536113981903  = 854.0
"1101011000",-- (0010010101) = 149.0     || 856.1938687102977  = 856.0
"1101011001",-- (0010010110) = 150.0     || 857.7228424532881  = 857.0
"1101011011",-- (0010010111) = 151.0     || 859.2405657145039  = 859.0
"1101011100",-- (0010011000) = 152.0     || 860.7470724321108  = 860.0
"1101011110",-- (0010011001) = 153.0     || 862.2423973763811  = 862.0
"1101011111",-- (0010011010) = 154.0     || 863.7265761310637  = 863.0
"1101100001",-- (0010011011) = 155.0     || 865.1996450748483  = 865.0
"1101100010",-- (0010011100) = 156.0     || 866.6616413629229  = 866.0
"1101100100",-- (0010011101) = 157.0     || 868.1126029086386  = 868.0
"1101100101",-- (0010011110) = 158.0     || 869.552568365279   = 869.0
"1101100110",-- (0010011111) = 159.0     || 870.9815771079438  = 870.0
"1101101000",-- (0010100000) = 160.0     || 872.39966921555    = 872.0
"1101101001",-- (0010100001) = 161.0     || 873.8068854529546  = 873.0
"1101101011",-- (0010100010) = 162.0     || 875.2032672532047  = 875.0
"1101101100",-- (0010100011) = 163.0     || 876.5888566999175  = 876.0
"1101101101",-- (0010100100) = 164.0     || 877.9636965097958  = 877.0
"1101101111",-- (0010100101) = 165.0     || 879.3278300152823  = 879.0
"1101110000",-- (0010100110) = 166.0     || 880.6813011473562  = 880.0
"1101110010",-- (0010100111) = 167.0     || 882.0241544184755  = 882.0
"1101110011",-- (0010101000) = 168.0     || 883.3564349056704  = 883.0
"1101110100",-- (0010101001) = 169.0     || 884.6781882337876  = 884.0
"1101110101",-- (0010101010) = 170.0     || 885.9894605588923  = 885.0
"1101110111",-- (0010101011) = 171.0     || 887.2902985518275  = 887.0
"1101111000",-- (0010101100) = 172.0     || 888.5807493819368  = 888.0
"1101111001",-- (0010101101) = 173.0     || 889.8608607009502  = 889.0
"1101111011",-- (0010101110) = 174.0     || 891.1306806270377  = 891.0
"1101111100",-- (0010101111) = 175.0     || 892.3902577290311  = 892.0
"1101111101",-- (0010110000) = 176.0     || 893.6396410108193  = 893.0
"1101111110",-- (0010110001) = 177.0     || 894.8788798959157  = 894.0
"1110000000",-- (0010110010) = 178.0     || 896.1080242122008  = 896.0
"1110000001",-- (0010110011) = 179.0     || 897.3271241768446  = 897.0
"1110000010",-- (0010110100) = 180.0     || 898.5362303814048  = 898.0
"1110000011",-- (0010110101) = 181.0     || 899.7353937771096  = 899.0
"1110000100",-- (0010110110) = 182.0     || 900.9246656603187  = 900.0
"1110000110",-- (0010110111) = 183.0     || 902.1040976581702  = 902.0
"1110000111",-- (0010111000) = 184.0     || 903.2737417144124  = 903.0
"1110001000",-- (0010111001) = 185.0     || 904.4336500754195  = 904.0
"1110001001",-- (0010111010) = 186.0     || 905.5838752763952  = 905.0
"1110001010",-- (0010111011) = 187.0     || 906.7244701277646  = 906.0
"1110001011",-- (0010111100) = 188.0     || 907.8554877017517  = 907.0
"1110001100",-- (0010111101) = 189.0     || 908.9769813191493  = 908.0
"1110001110",-- (0010111110) = 190.0     || 910.089004536276   = 910.0
"1110001111",-- (0010111111) = 191.0     || 911.1916111321227  = 911.0
"1110010000",-- (0011000000) = 192.0     || 912.2848550956924  = 912.0
"1110010001",-- (0011000001) = 193.0     || 913.3687906135259  = 913.0
"1110010010",-- (0011000010) = 194.0     || 914.4434720574222  = 914.0
"1110010011",-- (0011000011) = 195.0     || 915.5089539723472  = 915.0
"1110010100",-- (0011000100) = 196.0     || 916.5652910645325  = 916.0
"1110010101",-- (0011000101) = 197.0     || 917.6125381897674  = 917.0
"1110010110",-- (0011000110) = 198.0     || 918.6507503418776  = 918.0
"1110010111",-- (0011000111) = 199.0     || 919.6799826413957  = 919.0
"1110011000",-- (0011001000) = 200.0     || 920.7002903244222  = 920.0
"1110011001",-- (0011001001) = 201.0     || 921.7117287316719  = 921.0
"1110011010",-- (0011001010) = 202.0     || 922.7143532977135  = 922.0
"1110011011",-- (0011001011) = 203.0     || 923.7082195403926  = 923.0
"1110011100",-- (0011001100) = 204.0     || 924.6933830504461  = 924.0
"1110011101",-- (0011001101) = 205.0     || 925.6698994812991  = 925.0
"1110011110",-- (0011001110) = 206.0     || 926.6378245390507  = 926.0
"1110011111",-- (0011001111) = 207.0     || 927.5972139726426  = 927.0
"1110100000",-- (0011010000) = 208.0     || 928.5481235642126  = 928.0
"1110100001",-- (0011010001) = 209.0     || 929.4906091196307  = 929.0
"1110100010",-- (0011010010) = 210.0     || 930.4247264592166  = 930.0
"1110100011",-- (0011010011) = 211.0     || 931.3505314086389  = 931.0
"1110100100",-- (0011010100) = 212.0     || 932.2680797899932  = 932.0
"1110100101",-- (0011010101) = 213.0     || 933.1774274130588  = 933.0
"1110100110",-- (0011010110) = 214.0     || 934.0786300667327  = 934.0
"1110100110",-- (0011010111) = 215.0     || 934.9717435106389  = 934.0
"1110100111",-- (0011011000) = 216.0     || 935.856823466914   = 935.0
"1110101000",-- (0011011001) = 217.0     || 936.7339256121631  = 936.0
"1110101001",-- (0011011010) = 218.0     || 937.6031055695909  = 937.0
"1110101010",-- (0011011011) = 219.0     || 938.4644189012998  = 938.0
"1110101011",-- (0011011100) = 220.0     || 939.3179211007603  = 939.0
"1110101100",-- (0011011101) = 221.0     || 940.1636675854447  = 940.0
"1110101101",-- (0011011110) = 222.0     || 941.0017136896315  = 941.0
"1110101101",-- (0011011111) = 223.0     || 941.8321146573692  = 941.0
"1110101110",-- (0011100000) = 224.0     || 942.6549256356061  = 942.0
"1110101111",-- (0011100001) = 225.0     || 943.4702016674801  = 943.0
"1110110000",-- (0011100010) = 226.0     || 944.2779976857671  = 944.0
"1110110001",-- (0011100011) = 227.0     || 945.0783685064886  = 945.0
"1110110001",-- (0011100100) = 228.0     || 945.871368822674   = 945.0
"1110110010",-- (0011100101) = 229.0     || 946.657053198277   = 946.0
"1110110011",-- (0011100110) = 230.0     || 947.4354760622476  = 947.0
"1110110100",-- (0011100111) = 231.0     || 948.2066917027494  = 948.0
"1110110100",-- (0011101000) = 232.0     || 948.9707542615319  = 948.0
"1110110101",-- (0011101001) = 233.0     || 949.7277177284452  = 949.0
"1110110110",-- (0011101010) = 234.0     || 950.477635936104   = 950.0
"1110110111",-- (0011101011) = 235.0     || 951.2205625546922  = 951.0
"1110110111",-- (0011101100) = 236.0     || 951.9565510869112  = 951.0
"1110111000",-- (0011101101) = 237.0     || 952.6856548630682  = 952.0
"1110111001",-- (0011101110) = 238.0     || 953.4079270363015  = 953.0
"1110111010",-- (0011101111) = 239.0     || 954.1234205779442  = 954.0
"1110111010",-- (0011110000) = 240.0     || 954.8321882730198  = 954.0
"1110111011",-- (0011110001) = 241.0     || 955.5342827158725  = 955.0
"1110111100",-- (0011110010) = 242.0     || 956.229756305928   = 956.0
"1110111100",-- (0011110011) = 243.0     || 956.9186612435838  = 956.0
"1110111101",-- (0011110100) = 244.0     || 957.6010495262242  = 957.0
"1110111110",-- (0011110101) = 245.0     || 958.2769729443637  = 958.0
"1110111110",-- (0011110110) = 246.0     || 958.9464830779131  = 958.0
"1110111111",-- (0011110111) = 247.0     || 959.6096312925649  = 959.0
"1111000000",-- (0011111000) = 248.0     || 960.2664687363018  = 960.0
"1111000000",-- (0011111001) = 249.0     || 960.9170463360214  = 960.0
"1111000001",-- (0011111010) = 250.0     || 961.5614147942761  = 961.0
"1111000010",-- (0011111011) = 251.0     || 962.19962458613    = 962.0
"1111000010",-- (0011111100) = 252.0     || 962.831725956126   = 962.0
"1111000011",-- (0011111101) = 253.0     || 963.4577689153637  = 963.0
"1111000100",-- (0011111110) = 254.0     || 964.0778032386867  = 964.0
"1111000100",-- (0011111111) = 255.0     || 964.6918784619783  = 964.0
"1111000101",-- (0100000000) = 256.0     || 965.3000438795584  = 965.0
"1111000101",-- (0100000001) = 257.0     || 965.902348541689   = 965.0
"1111000110",-- (0100000010) = 258.0     || 966.4988412521765  = 966.0
"1111000111",-- (0100000011) = 259.0     || 967.089570566078   = 967.0
"1111000111",-- (0100000100) = 260.0     || 967.674584787503   = 967.0
"1111001000",-- (0100000101) = 261.0     || 968.2539319675117  = 968.0
"1111001000",-- (0100000110) = 262.0     || 968.8276599021106  = 968.0
"1111001001",-- (0100000111) = 263.0     || 969.395816130337   = 969.0
"1111001001",-- (0100001000) = 264.0     || 969.9584479324386  = 969.0
"1111001010",-- (0100001001) = 265.0     || 970.5156023281401  = 970.0
"1111001011",-- (0100001010) = 266.0     || 971.067326074998   = 971.0
"1111001011",-- (0100001011) = 267.0     || 971.6136656668439  = 971.0
"1111001100",-- (0100001100) = 268.0     || 972.1546673323082  = 972.0
"1111001100",-- (0100001101) = 269.0     || 972.6903770334309  = 972.0
"1111001101",-- (0100001110) = 270.0     || 973.2208404643516  = 973.0
"1111001101",-- (0100001111) = 271.0     || 973.7461030500784  = 973.0
"1111001110",-- (0100010000) = 272.0     || 974.2662099453377  = 974.0
"1111001110",-- (0100010001) = 273.0     || 974.7812060334975  = 974.0
"1111001111",-- (0100010010) = 274.0     || 975.2911359255671  = 975.0
"1111001111",-- (0100010011) = 275.0     || 975.7960439592713  = 975.0
"1111010000",-- (0100010100) = 276.0     || 976.2959741981939  = 976.0
"1111010000",-- (0100010101) = 277.0     || 976.7909704309935  = 976.0
"1111010001",-- (0100010110) = 278.0     || 977.2810761706882  = 977.0
"1111010001",-- (0100010111) = 279.0     || 977.7663346540068  = 977.0
"1111010010",-- (0100011000) = 280.0     || 978.2467888408062  = 978.0
"1111010010",-- (0100011001) = 281.0     || 978.7224814135537  = 978.0
"1111010011",-- (0100011010) = 282.0     || 979.1934547768728  = 979.0
"1111010011",-- (0100011011) = 283.0     || 979.6597510571488  = 979.0
"1111010100",-- (0100011100) = 284.0     || 980.121412102197   = 980.0
"1111010100",-- (0100011101) = 285.0     || 980.578479480989   = 980.0
"1111010101",-- (0100011110) = 286.0     || 981.0309944834348  = 981.0
"1111010101",-- (0100011111) = 287.0     || 981.4789981202252  = 981.0
"1111010101",-- (0100100000) = 288.0     || 981.9225311227239  = 981.0
"1111010110",-- (0100100001) = 289.0     || 982.3616339429177  = 982.0
"1111010110",-- (0100100010) = 290.0     || 982.7963467534173  = 982.0
"1111010111",-- (0100100011) = 291.0     || 983.2267094475075  = 983.0
"1111010111",-- (0100100100) = 292.0     || 983.6527616392508  = 983.0
"1111011000",-- (0100100101) = 293.0     || 984.0745426636364  = 984.0
"1111011000",-- (0100100110) = 294.0     || 984.4920915767773  = 984.0
"1111011000",-- (0100100111) = 295.0     || 984.905447156156   = 984.0
"1111011001",-- (0100101000) = 296.0     || 985.3146479009108  = 985.0
"1111011001",-- (0100101001) = 297.0     || 985.7197320321698  = 985.0
"1111011010",-- (0100101010) = 298.0     || 986.1207374934262  = 986.0
"1111011010",-- (0100101011) = 299.0     || 986.5177019509538  = 986.0
"1111011010",-- (0100101100) = 300.0     || 986.9106627942659  = 986.0
"1111011011",-- (0100101101) = 301.0     || 987.2996571366103  = 987.0
"1111011011",-- (0100101110) = 302.0     || 987.6847218155059  = 987.0
"1111011100",-- (0100101111) = 303.0     || 988.0658933933124  = 988.0
"1111011100",-- (0100110000) = 304.0     || 988.4432081578418  = 988.0
"1111011100",-- (0100110001) = 305.0     || 988.8167021229988  = 988.0
"1111011101",-- (0100110010) = 306.0     || 989.18641102946    = 989.0
"1111011101",-- (0100110011) = 307.0     || 989.5523703453848  = 989.0
"1111011101",-- (0100110100) = 308.0     || 989.9146152671578  = 989.0
"1111011110",-- (0100110101) = 309.0     || 990.2731807201634  = 990.0
"1111011110",-- (0100110110) = 310.0     || 990.62810135959    = 990.0
"1111011110",-- (0100110111) = 311.0     || 990.9794115712646  = 990.0
"1111011111",-- (0100111000) = 312.0     || 991.3271454725144  = 991.0
"1111011111",-- (0100111001) = 313.0     || 991.6713369130579  = 991.0
"1111100000",-- (0100111010) = 314.0     || 992.0120194759197  = 992.0
"1111100000",-- (0100111011) = 315.0     || 992.3492264783757  = 992.0
"1111100000",-- (0100111100) = 316.0     || 992.6829909729187  = 992.0
"1111100001",-- (0100111101) = 317.0     || 993.0133457482501  = 993.0
"1111100001",-- (0100111110) = 318.0     || 993.3403233302969  = 993.0
"1111100001",-- (0100111111) = 319.0     || 993.6639559832472  = 993.0
"1111100001",-- (0101000000) = 320.0     || 993.9842757106111  = 993.0
"1111100010",-- (0101000001) = 321.0     || 994.3013142563004  = 994.0
"1111100010",-- (0101000010) = 322.0     || 994.6151031057299  = 994.0
"1111100010",-- (0101000011) = 323.0     || 994.9256734869374  = 994.0
"1111100011",-- (0101000100) = 324.0     || 995.2330563717226  = 995.0
"1111100011",-- (0101000101) = 325.0     || 995.537282476805   = 995.0
"1111100011",-- (0101000110) = 326.0     || 995.8383822649976  = 995.0
"1111100100",-- (0101000111) = 327.0     || 996.1363859463987  = 996.0
"1111100100",-- (0101001000) = 328.0     || 996.4313234795991  = 996.0
"1111100100",-- (0101001001) = 329.0     || 996.7232245729043  = 996.0
"1111100101",-- (0101001010) = 330.0     || 997.0121186855732  = 997.0
"1111100101",-- (0101001011) = 331.0     || 997.2980350290688  = 997.0
"1111100101",-- (0101001100) = 332.0     || 997.5810025683228  = 997.0
"1111100101",-- (0101001101) = 333.0     || 997.8610500230146  = 997.0
"1111100110",-- (0101001110) = 334.0     || 998.138205868861   = 998.0
"1111100110",-- (0101001111) = 335.0     || 998.4124983389181  = 998.0
"1111100110",-- (0101010000) = 336.0     || 998.6839554248953  = 998.0
"1111100110",-- (0101010001) = 337.0     || 998.9526048784782  = 998.0
"1111100111",-- (0101010010) = 338.0     || 999.2184742126626  = 999.0
"1111100111",-- (0101010011) = 339.0     || 999.4815907030982  = 999.0
"1111100111",-- (0101010100) = 340.0     || 999.7419813894406  = 999.0
"1111100111",-- (0101010101) = 341.0     || 999.999673076713   = 999.0
"1111101000",-- (0101010110) = 342.0     || 1000.2546923366741 = 1000.0
"1111101000",-- (0101010111) = 343.0     || 1000.5070655091959 = 1000.0
"1111101000",-- (0101011000) = 344.0     || 1000.7568187036459 = 1000.0
"1111101001",-- (0101011001) = 345.0     || 1001.0039778002779 = 1001.0
"1111101001",-- (0101011010) = 346.0     || 1001.2485684516289 = 1001.0
"1111101001",-- (0101011011) = 347.0     || 1001.49061608392   = 1001.0
"1111101001",-- (0101011100) = 348.0     || 1001.7301458984648 = 1001.0
"1111101001",-- (0101011101) = 349.0     || 1001.9671828730807 = 1001.0
"1111101010",-- (0101011110) = 350.0     || 1002.2017517635061 = 1002.0
"1111101010",-- (0101011111) = 351.0     || 1002.433877104821  = 1002.0
"1111101010",-- (0101100000) = 352.0     || 1002.6635832128712 = 1002.0
"1111101010",-- (0101100001) = 353.0     || 1002.8908941856961 = 1002.0
"1111101011",-- (0101100010) = 354.0     || 1003.1158339049592 = 1003.0
"1111101011",-- (0101100011) = 355.0     || 1003.3384260373812 = 1003.0
"1111101011",-- (0101100100) = 356.0     || 1003.558694036175  = 1003.0
"1111101011",-- (0101100101) = 357.0     || 1003.7766611424836 = 1003.0
"1111101011",-- (0101100110) = 358.0     || 1003.9923503868179 = 1003.0
"1111101100",-- (0101100111) = 359.0     || 1004.2057845904972 = 1004.0
"1111101100",-- (0101101000) = 360.0     || 1004.4169863670899 = 1004.0
"1111101100",-- (0101101001) = 361.0     || 1004.6259781238534 = 1004.0
"1111101100",-- (0101101010) = 362.0     || 1004.8327820631783 = 1004.0
"1111101101",-- (0101101011) = 363.0     || 1005.0374201840277 = 1005.0
"1111101101",-- (0101101100) = 364.0     || 1005.2399142833789 = 1005.0
"1111101101",-- (0101101101) = 365.0     || 1005.4402859576641 = 1005.0
"1111101101",-- (0101101110) = 366.0     || 1005.6385566042106 = 1005.0
"1111101101",-- (0101101111) = 367.0     || 1005.8347474226789 = 1005.0
"1111101110",-- (0101110000) = 368.0     || 1006.0288794164999 = 1006.0
"1111101110",-- (0101110001) = 369.0     || 1006.22097339431   = 1006.0
"1111101110",-- (0101110010) = 370.0     || 1006.4110499713861 = 1006.0
"1111101110",-- (0101110011) = 371.0     || 1006.5991295710755 = 1006.0
"1111101110",-- (0101110100) = 372.0     || 1006.7852324262268 = 1006.0
"1111101110",-- (0101110101) = 373.0     || 1006.9693785806155 = 1006.0
"1111101111",-- (0101110110) = 374.0     || 1007.1515878903675 = 1007.0
"1111101111",-- (0101110111) = 375.0     || 1007.3318800253813 = 1007.0
"1111101111",-- (0101111000) = 376.0     || 1007.510274470745  = 1007.0
"1111101111",-- (0101111001) = 377.0     || 1007.6867905281505 = 1007.0
"1111101111",-- (0101111010) = 378.0     || 1007.861447317304  = 1007.0
"1111110000",-- (0101111011) = 379.0     || 1008.0342637773346 = 1008.0
"1111110000",-- (0101111100) = 380.0     || 1008.2052586681946 = 1008.0
"1111110000",-- (0101111101) = 381.0     || 1008.3744505720617 = 1008.0
"1111110000",-- (0101111110) = 382.0     || 1008.5418578947312 = 1008.0
"1111110000",-- (0101111111) = 383.0     || 1008.7074988670073 = 1008.0
"1111110000",-- (0110000000) = 384.0     || 1008.8713915460884 = 1008.0
"1111110001",-- (0110000001) = 385.0     || 1009.0335538169488 = 1009.0
"1111110001",-- (0110000010) = 386.0     || 1009.1940033937138 = 1009.0
"1111110001",-- (0110000011) = 387.0     || 1009.3527578210313 = 1009.0
"1111110001",-- (0110000100) = 388.0     || 1009.509834475438  = 1009.0
"1111110001",-- (0110000101) = 389.0     || 1009.6652505667183 = 1009.0
"1111110001",-- (0110000110) = 390.0     || 1009.8190231392618 = 1009.0
"1111110001",-- (0110000111) = 391.0     || 1009.9711690734117 = 1009.0
"1111110010",-- (0110001000) = 392.0     || 1010.1217050868082 = 1010.0
"1111110010",-- (0110001001) = 393.0     || 1010.2706477357281 = 1010.0
"1111110010",-- (0110001010) = 394.0     || 1010.4180134164163 = 1010.0
"1111110010",-- (0110001011) = 395.0     || 1010.5638183664117 = 1010.0
"1111110010",-- (0110001100) = 396.0     || 1010.7080786658692 = 1010.0
"1111110010",-- (0110001101) = 397.0     || 1010.8508102388718 = 1010.0
"1111110010",-- (0110001110) = 398.0     || 1010.9920288547396 = 1010.0
"1111110011",-- (0110001111) = 399.0     || 1011.1317501293308 = 1011.0
"1111110011",-- (0110010000) = 400.0     || 1011.2699895263377 = 1011.0
"1111110011",-- (0110010001) = 401.0     || 1011.4067623585738 = 1011.0
"1111110011",-- (0110010010) = 402.0     || 1011.5420837892569 = 1011.0
"1111110011",-- (0110010011) = 403.0     || 1011.6759688332836 = 1011.0
"1111110011",-- (0110010100) = 404.0     || 1011.8084323584985 = 1011.0
"1111110011",-- (0110010101) = 405.0     || 1011.9394890869559 = 1011.0
"1111110100",-- (0110010110) = 406.0     || 1012.0691535961739 = 1012.0
"1111110100",-- (0110010111) = 407.0     || 1012.1974403203832 = 1012.0
"1111110100",-- (0110011000) = 408.0     || 1012.3243635517679 = 1012.0
"1111110100",-- (0110011001) = 409.0     || 1012.449937441699  = 1012.0
"1111110100",-- (0110011010) = 410.0     || 1012.574176001962  = 1012.0
"1111110100",-- (0110011011) = 411.0     || 1012.6970931059757 = 1012.0
"1111110100",-- (0110011100) = 412.0     || 1012.8187024900059 = 1012.0
"1111110100",-- (0110011101) = 413.0     || 1012.9390177543694 = 1012.0
"1111110101",-- (0110011110) = 414.0     || 1013.0580523646333 = 1013.0
"1111110101",-- (0110011111) = 415.0     || 1013.175819652805  = 1013.0
"1111110101",-- (0110100000) = 416.0     || 1013.2923328185158 = 1013.0
"1111110101",-- (0110100001) = 417.0     || 1013.4076049301974 = 1013.0
"1111110101",-- (0110100010) = 418.0     || 1013.5216489262497 = 1013.0
"1111110101",-- (0110100011) = 419.0     || 1013.6344776162026 = 1013.0
"1111110101",-- (0110100100) = 420.0     || 1013.7461036818706 = 1013.0
"1111110101",-- (0110100101) = 421.0     || 1013.8565396784979 = 1013.0
"1111110101",-- (0110100110) = 422.0     || 1013.9657980358976 = 1013.0
"1111110110",-- (0110100111) = 423.0     || 1014.0738910595833 = 1014.0
"1111110110",-- (0110101000) = 424.0     || 1014.1808309318931 = 1014.0
"1111110110",-- (0110101001) = 425.0     || 1014.2866297131056 = 1014.0
"1111110110",-- (0110101010) = 426.0     || 1014.3912993425492 = 1014.0
"1111110110",-- (0110101011) = 427.0     || 1014.4948516397022 = 1014.0
"1111110110",-- (0110101100) = 428.0     || 1014.5972983052877 = 1014.0
"1111110110",-- (0110101101) = 429.0     || 1014.698650922359  = 1014.0
"1111110110",-- (0110101110) = 430.0     || 1014.7989209573784 = 1014.0
"1111110110",-- (0110101111) = 431.0     || 1014.898119761288  = 1014.0
"1111110110",-- (0110110000) = 432.0     || 1014.9962585705729 = 1014.0
"1111110111",-- (0110110001) = 433.0     || 1015.0933485083176 = 1015.0
"1111110111",-- (0110110010) = 434.0     || 1015.1894005852535 = 1015.0
"1111110111",-- (0110110011) = 435.0     || 1015.2844257007999 = 1015.0
"1111110111",-- (0110110100) = 436.0     || 1015.3784346440973 = 1015.0
"1111110111",-- (0110110101) = 437.0     || 1015.471438095032  = 1015.0
"1111110111",-- (0110110110) = 438.0     || 1015.5634466252556 = 1015.0
"1111110111",-- (0110110111) = 439.0     || 1015.6544706991936 = 1015.0
"1111110111",-- (0110111000) = 440.0     || 1015.7445206750499 = 1015.0
"1111110111",-- (0110111001) = 441.0     || 1015.8336068058012 = 1015.0
"1111110111",-- (0110111010) = 442.0     || 1015.9217392401853 = 1015.0
"1111111000",-- (0110111011) = 443.0     || 1016.0089280236809 = 1016.0
"1111111000",-- (0110111100) = 444.0     || 1016.095183099482  = 1016.0
"1111111000",-- (0110111101) = 445.0     || 1016.1805143094608 = 1016.0
"1111111000",-- (0110111110) = 446.0     || 1016.2649313951282 = 1016.0
"1111111000",-- (0110111111) = 447.0     || 1016.348443998583  = 1016.0
"1111111000",-- (0111000000) = 448.0     || 1016.4310616634554 = 1016.0
"1111111000",-- (0111000001) = 449.0     || 1016.5127938358424 = 1016.0
"1111111000",-- (0111000010) = 450.0     || 1016.5936498652375 = 1016.0
"1111111000",-- (0111000011) = 451.0     || 1016.6736390054499 = 1016.0
"1111111000",-- (0111000100) = 452.0     || 1016.7527704155198 = 1016.0
"1111111000",-- (0111000101) = 453.0     || 1016.831053160624  = 1016.0
"1111111000",-- (0111000110) = 454.0     || 1016.9084962129755 = 1016.0
"1111111000",-- (0111000111) = 455.0     || 1016.9851084527155 = 1016.0
"1111111001",-- (0111001000) = 456.0     || 1017.0608986687981 = 1017.0
"1111111001",-- (0111001001) = 457.0     || 1017.1358755598674 = 1017.0
"1111111001",-- (0111001010) = 458.0     || 1017.2100477351283 = 1017.0
"1111111001",-- (0111001011) = 459.0     || 1017.2834237152106 = 1017.0
"1111111001",-- (0111001100) = 460.0     || 1017.3560119330236 = 1017.0
"1111111001",-- (0111001101) = 461.0     || 1017.4278207346058 = 1017.0
"1111111001",-- (0111001110) = 462.0     || 1017.4988583799682 = 1017.0
"1111111001",-- (0111001111) = 463.0     || 1017.5691330439271 = 1017.0
"1111111001",-- (0111010000) = 464.0     || 1017.6386528169342 = 1017.0
"1111111001",-- (0111010001) = 465.0     || 1017.7074257058968 = 1017.0
"1111111001",-- (0111010010) = 466.0     || 1017.7754596349921 = 1017.0
"1111111001",-- (0111010011) = 467.0     || 1017.842762446475  = 1017.0
"1111111001",-- (0111010100) = 468.0     || 1017.9093419014779 = 1017.0
"1111111001",-- (0111010101) = 469.0     || 1017.9752056808048 = 1017.0
"1111111010",-- (0111010110) = 470.0     || 1018.0403613857188 = 1018.0
"1111111010",-- (0111010111) = 471.0     || 1018.1048165387213 = 1018.0
"1111111010",-- (0111011000) = 472.0     || 1018.1685785843259 = 1018.0
"1111111010",-- (0111011001) = 473.0     || 1018.231654889826  = 1018.0
"1111111010",-- (0111011010) = 474.0     || 1018.2940527460535 = 1018.0
"1111111010",-- (0111011011) = 475.0     || 1018.3557793681337 = 1018.0
"1111111010",-- (0111011100) = 476.0     || 1018.4168418962317 = 1018.0
"1111111010",-- (0111011101) = 477.0     || 1018.4772473962934 = 1018.0
"1111111010",-- (0111011110) = 478.0     || 1018.537002860779  = 1018.0
"1111111010",-- (0111011111) = 479.0     || 1018.5961152093912 = 1018.0
"1111111010",-- (0111100000) = 480.0     || 1018.6545912897963 = 1018.0
"1111111010",-- (0111100001) = 481.0     || 1018.7124378783382 = 1018.0
"1111111010",-- (0111100010) = 482.0     || 1018.7696616807478 = 1018.0
"1111111010",-- (0111100011) = 483.0     || 1018.826269332846  = 1018.0
"1111111010",-- (0111100100) = 484.0     || 1018.8822674012375 = 1018.0
"1111111010",-- (0111100101) = 485.0     || 1018.9376623840026 = 1018.0
"1111111010",-- (0111100110) = 486.0     || 1018.9924607113792 = 1018.0
"1111111011",-- (0111100111) = 487.0     || 1019.0466687464418 = 1019.0
"1111111011",-- (0111101000) = 488.0     || 1019.100292785772  = 1019.0
"1111111011",-- (0111101001) = 489.0     || 1019.1533390601235 = 1019.0
"1111111011",-- (0111101010) = 490.0     || 1019.2058137350822 = 1019.0
"1111111011",-- (0111101011) = 491.0     || 1019.2577229117193 = 1019.0
"1111111011",-- (0111101100) = 492.0     || 1019.3090726272382 = 1019.0
"1111111011",-- (0111101101) = 493.0     || 1019.3598688556164 = 1019.0
"1111111011",-- (0111101110) = 494.0     || 1019.4101175082418 = 1019.0
"1111111011",-- (0111101111) = 495.0     || 1019.4598244345409 = 1019.0
"1111111011",-- (0111110000) = 496.0     || 1019.5089954226046 = 1019.0
"1111111011",-- (0111110001) = 497.0     || 1019.5576361998055 = 1019.0
"1111111011",-- (0111110010) = 498.0     || 1019.6057524334109 = 1019.0
"1111111011",-- (0111110011) = 499.0     || 1019.6533497311892 = 1019.0
"1111111011",-- (0111110100) = 500.0     || 1019.7004336420127 = 1019.0
"1111111011",-- (0111110101) = 501.0     || 1019.747009656452  = 1019.0
"1111111011",-- (0111110110) = 502.0     || 1019.7930832073665 = 1019.0
"1111111011",-- (0111110111) = 503.0     || 1019.83865967049   = 1019.0
"1111111011",-- (0111111000) = 504.0     || 1019.8837443650087 = 1019.0
"1111111011",-- (0111111001) = 505.0     || 1019.9283425541373 = 1019.0
"1111111011",-- (0111111010) = 506.0     || 1019.9724594456846 = 1019.0
"1111111100",-- (0111111011) = 507.0     || 1020.0161001926191 = 1020.0
"1111111100",-- (0111111100) = 508.0     || 1020.0592698936263 = 1020.0
"1111111100",-- (0111111101) = 509.0     || 1020.1019735936605 = 1020.0
"1111111100",-- (0111111110) = 510.0     || 1020.144216284494  = 1020.0
"1111111100",-- (0111111111) = 511.0     || 1020.1860029052572 = 1020.0
"0000000011",-- (1000000000) = -512.0    || 3.7726616570224527 = 3.0
"0000000011",-- (1000000001) = -511.0    || 3.813997094742907  = 3.0
"0000000011",-- (1000000010) = -510.0    || 3.855783715506047  = 3.0
"0000000011",-- (1000000011) = -509.0    || 3.8980264063393055 = 3.0
"0000000011",-- (1000000100) = -508.0    || 3.9407301063736497 = 3.0
"0000000011",-- (1000000101) = -507.0    || 3.9838998073807748 = 3.0
"0000000100",-- (1000000110) = -506.0    || 4.027540554315391  = 4.0
"0000000100",-- (1000000111) = -505.0    || 4.071657445862708  = 4.0
"0000000100",-- (1000001000) = -504.0    || 4.11625563499111   = 4.0
"0000000100",-- (1000001001) = -503.0    || 4.1613403295100895 = 4.0
"0000000100",-- (1000001010) = -502.0    || 4.20691679263348   = 4.0
"0000000100",-- (1000001011) = -501.0    || 4.252990343548004  = 4.0
"0000000100",-- (1000001100) = -500.0    || 4.299566357987193  = 4.0
"0000000100",-- (1000001101) = -499.0    || 4.346650268810732  = 4.0
"0000000100",-- (1000001110) = -498.0    || 4.394247566589228  = 4.0
"0000000100",-- (1000001111) = -497.0    || 4.442363800194505  = 4.0
"0000000100",-- (1000010000) = -496.0    || 4.491004577395397  = 4.0
"0000000100",-- (1000010001) = -495.0    || 4.54017556545913   = 4.0
"0000000100",-- (1000010010) = -494.0    || 4.58988249175832   = 4.0
"0000000100",-- (1000010011) = -493.0    || 4.640131144383588  = 4.0
"0000000100",-- (1000010100) = -492.0    || 4.690927372761929  = 4.0
"0000000100",-- (1000010101) = -491.0    || 4.7422770882807574 = 4.0
"0000000100",-- (1000010110) = -490.0    || 4.794186264917747  = 4.0
"0000000100",-- (1000010111) = -489.0    || 4.846660939876494  = 4.0
"0000000100",-- (1000011000) = -488.0    || 4.899707214228002  = 4.0
"0000000100",-- (1000011001) = -487.0    || 4.953331253558106  = 4.0
"0000000101",-- (1000011010) = -486.0    || 5.00753928862079   = 5.0
"0000000101",-- (1000011011) = -485.0    || 5.0623376159974915 = 5.0
"0000000101",-- (1000011100) = -484.0    || 5.1177325987624345 = 5.0
"0000000101",-- (1000011101) = -483.0    || 5.173730667153973  = 5.0
"0000000101",-- (1000011110) = -482.0    || 5.230338319252091  = 5.0
"0000000101",-- (1000011111) = -481.0    || 5.287562121661977  = 5.0
"0000000101",-- (1000100000) = -480.0    || 5.345408710203799  = 5.0
"0000000101",-- (1000100001) = -479.0    || 5.403884790608691  = 5.0
"0000000101",-- (1000100010) = -478.0    || 5.462997139220963  = 5.0
"0000000101",-- (1000100011) = -477.0    || 5.5227526037066506 = 5.0
"0000000101",-- (1000100100) = -476.0    || 5.583158103768338  = 5.0
"0000000101",-- (1000100101) = -475.0    || 5.6442206318663874 = 5.0
"0000000101",-- (1000100110) = -474.0    || 5.705947253946553  = 5.0
"0000000101",-- (1000100111) = -473.0    || 5.768345110174028  = 5.0
"0000000101",-- (1000101000) = -472.0    || 5.831421415674016  = 5.0
"0000000101",-- (1000101001) = -471.0    || 5.895183461278771  = 5.0
"0000000101",-- (1000101010) = -470.0    || 5.959638614281224  = 5.0
"0000000110",-- (1000101011) = -469.0    || 6.024794319195192  = 6.0
"0000000110",-- (1000101100) = -468.0    || 6.090658098522197  = 6.0
"0000000110",-- (1000101101) = -467.0    || 6.1572375535250075 = 6.0
"0000000110",-- (1000101110) = -466.0    || 6.224540365007817  = 6.0
"0000000110",-- (1000101111) = -465.0    || 6.292574294103197  = 6.0
"0000000110",-- (1000110000) = -464.0    || 6.36134718306582   = 6.0
"0000000110",-- (1000110001) = -463.0    || 6.4308669560729586 = 6.0
"0000000110",-- (1000110010) = -462.0    || 6.501141620031886  = 6.0
"0000000110",-- (1000110011) = -461.0    || 6.572179265394097  = 6.0
"0000000110",-- (1000110100) = -460.0    || 6.6439880669764655 = 6.0
"0000000110",-- (1000110101) = -459.0    || 6.716576284789339  = 6.0
"0000000110",-- (1000110110) = -458.0    || 6.789952264871589  = 6.0
"0000000110",-- (1000110111) = -457.0    || 6.864124440132721  = 6.0
"0000000110",-- (1000111000) = -456.0    || 6.93910133120196   = 6.0
"0000000111",-- (1000111001) = -455.0    || 7.0148915472844475 = 7.0
"0000000111",-- (1000111010) = -454.0    || 7.09150378702452   = 7.0
"0000000111",-- (1000111011) = -453.0    || 7.168946839376097  = 7.0
"0000000111",-- (1000111100) = -452.0    || 7.247229584480292  = 7.0
"0000000111",-- (1000111101) = -451.0    || 7.326360994550133  = 7.0
"0000000111",-- (1000111110) = -450.0    || 7.406350134762546  = 7.0
"0000000111",-- (1000111111) = -449.0    || 7.4872061641575565 = 7.0
"0000000111",-- (1001000000) = -448.0    || 7.568938336544744  = 7.0
"0000000111",-- (1001000001) = -447.0    || 7.651556001417048  = 7.0
"0000000111",-- (1001000010) = -446.0    || 7.735068604871815  = 7.0
"0000000111",-- (1001000011) = -445.0    || 7.819485690539225  = 7.0
"0000000111",-- (1001000100) = -444.0    || 7.904816900518086  = 7.0
"0000000111",-- (1001000101) = -443.0    || 7.991071976318964  = 7.0
"0000001000",-- (1001000110) = -442.0    || 8.078260759814793  = 8.0
"0000001000",-- (1001000111) = -441.0    || 8.166393194198843  = 8.0
"0000001000",-- (1001001000) = -440.0    || 8.25547932495016   = 8.0
"0000001000",-- (1001001001) = -439.0    || 8.345529300806469  = 8.0
"0000001000",-- (1001001010) = -438.0    || 8.436553374744511  = 8.0
"0000001000",-- (1001001011) = -437.0    || 8.528561904967964  = 8.0
"0000001000",-- (1001001100) = -436.0    || 8.621565355902773  = 8.0
"0000001000",-- (1001001101) = -435.0    || 8.715574299200053  = 8.0
"0000001000",-- (1001001110) = -434.0    || 8.810599414746521  = 8.0
"0000001000",-- (1001001111) = -433.0    || 8.906651491682428  = 8.0
"0000001001",-- (1001010000) = -432.0    || 9.003741429427121  = 9.0
"0000001001",-- (1001010001) = -431.0    || 9.10188023871209   = 9.0
"0000001001",-- (1001010010) = -430.0    || 9.201079042621618  = 9.0
"0000001001",-- (1001010011) = -429.0    || 9.301349077641005  = 9.0
"0000001001",-- (1001010100) = -428.0    || 9.402701694712315  = 9.0
"0000001001",-- (1001010101) = -427.0    || 9.5051483602978    = 9.0
"0000001001",-- (1001010110) = -426.0    || 9.608700657450804  = 9.0
"0000001001",-- (1001010111) = -425.0    || 9.71337028689429   = 9.0
"0000001001",-- (1001011000) = -424.0    || 9.819169068106948  = 9.0
"0000001001",-- (1001011001) = -423.0    || 9.926108940416805  = 9.0
"0000001010",-- (1001011010) = -422.0    || 10.034201964102516 = 10.0
"0000001010",-- (1001011011) = -421.0    || 10.143460321502106 = 10.0
"0000001010",-- (1001011100) = -420.0    || 10.253896318129293 = 10.0
"0000001010",-- (1001011101) = -419.0    || 10.365522383797353 = 10.0
"0000001010",-- (1001011110) = -418.0    || 10.478351073750474 = 10.0
"0000001010",-- (1001011111) = -417.0    || 10.592395069802668 = 10.0
"0000001010",-- (1001100000) = -416.0    || 10.707667181484105 = 10.0
"0000001010",-- (1001100001) = -415.0    || 10.824180347194954 = 10.0
"0000001010",-- (1001100010) = -414.0    || 10.941947635366658 = 10.0
"0000001011",-- (1001100011) = -413.0    || 11.06098224563058  = 11.0
"0000001011",-- (1001100100) = -412.0    || 11.181297509994149 = 11.0
"0000001011",-- (1001100101) = -411.0    || 11.302906894024261 = 11.0
"0000001011",-- (1001100110) = -410.0    || 11.425823998038052 = 11.0
"0000001011",-- (1001100111) = -409.0    || 11.550062558300981 = 11.0
"0000001011",-- (1001101000) = -408.0    || 11.675636448232122 = 11.0
"0000001011",-- (1001101001) = -407.0    || 11.802559679616763 = 11.0
"0000001011",-- (1001101010) = -406.0    || 11.9308464038261   = 11.0
"0000001100",-- (1001101011) = -405.0    || 12.060510913044094 = 12.0
"0000001100",-- (1001101100) = -404.0    || 12.191567641501429 = 12.0
"0000001100",-- (1001101101) = -403.0    || 12.324031166716452 = 12.0
"0000001100",-- (1001101110) = -402.0    || 12.457916210743189 = 12.0
"0000001100",-- (1001101111) = -401.0    || 12.593237641426189 = 12.0
"0000001100",-- (1001110000) = -400.0    || 12.73001047366228  = 12.0
"0000001100",-- (1001110001) = -399.0    || 12.86824987066913  = 12.0
"0000001101",-- (1001110010) = -398.0    || 13.007971145260496 = 13.0
"0000001101",-- (1001110011) = -397.0    || 13.149189761128218 = 13.0
"0000001101",-- (1001110100) = -396.0    || 13.291921334130743 = 13.0
"0000001101",-- (1001110101) = -395.0    || 13.43618163358818  = 13.0
"0000001101",-- (1001110110) = -394.0    || 13.581986583583808 = 13.0
"0000001101",-- (1001110111) = -393.0    || 13.729352264271883 = 13.0
"0000001101",-- (1001111000) = -392.0    || 13.878294913191807 = 13.0
"0000001110",-- (1001111001) = -391.0    || 14.02883092658837  = 14.0
"0000001110",-- (1001111010) = -390.0    || 14.180976860738124 = 14.0
"0000001110",-- (1001111011) = -389.0    || 14.334749433281733 = 14.0
"0000001110",-- (1001111100) = -388.0    || 14.490165524562121 = 14.0
"0000001110",-- (1001111101) = -387.0    || 14.647242178968547 = 14.0
"0000001110",-- (1001111110) = -386.0    || 14.805996606286167 = 14.0
"0000001110",-- (1001111111) = -385.0    || 14.966446183051216 = 14.0
"0000001111",-- (1010000000) = -384.0    || 15.128608453911621 = 15.0
"0000001111",-- (1010000001) = -383.0    || 15.292501132992799 = 15.0
"0000001111",-- (1010000010) = -382.0    || 15.458142105268783 = 15.0
"0000001111",-- (1010000011) = -381.0    || 15.62554942793822  = 15.0
"0000001111",-- (1010000100) = -380.0    || 15.794741331805325 = 15.0
"0000001111",-- (1010000101) = -379.0    || 15.965736222665566 = 15.0
"0000010000",-- (1010000110) = -378.0    || 16.138552682695934 = 16.0
"0000010000",-- (1010000111) = -377.0    || 16.313209471849596 = 16.0
"0000010000",-- (1010001000) = -376.0    || 16.489725529254947 = 16.0
"0000010000",-- (1010001001) = -375.0    || 16.668119974618623 = 16.0
"0000010000",-- (1010001010) = -374.0    || 16.848412109632523 = 16.0
"0000010001",-- (1010001011) = -373.0    || 17.030621419384605 = 17.0
"0000010001",-- (1010001100) = -372.0    || 17.21476757377313  = 17.0
"0000010001",-- (1010001101) = -371.0    || 17.40087042892449  = 17.0
"0000010001",-- (1010001110) = -370.0    || 17.588950028614047 = 17.0
"0000010001",-- (1010001111) = -369.0    || 17.779026605690017 = 17.0
"0000010001",-- (1010010000) = -368.0    || 17.971120583500173 = 17.0
"0000010010",-- (1010010001) = -367.0    || 18.16525257732098  = 18.0
"0000010010",-- (1010010010) = -366.0    || 18.361443395789284 = 18.0
"0000010010",-- (1010010011) = -365.0    || 18.559714042335898 = 18.0
"0000010010",-- (1010010100) = -364.0    || 18.76008571662118  = 18.0
"0000010010",-- (1010010101) = -363.0    || 18.962579815972237 = 18.0
"0000010011",-- (1010010110) = -362.0    || 19.16721793682152  = 19.0
"0000010011",-- (1010010111) = -361.0    || 19.374021876146482 = 19.0
"0000010011",-- (1010011000) = -360.0    || 19.583013632910248 = 19.0
"0000010011",-- (1010011001) = -359.0    || 19.7942154095027   = 19.0
"0000010100",-- (1010011010) = -358.0    || 20.007649613182075 = 20.0
"0000010100",-- (1010011011) = -357.0    || 20.223338857516453 = 20.0
"0000010100",-- (1010011100) = -356.0    || 20.441305963825027 = 20.0
"0000010100",-- (1010011101) = -355.0    || 20.66157396261888  = 20.0
"0000010100",-- (1010011110) = -354.0    || 20.88416609504077  = 20.0
"0000010101",-- (1010011111) = -353.0    || 21.10910581430384  = 21.0
"0000010101",-- (1010100000) = -352.0    || 21.336416787128762 = 21.0
"0000010101",-- (1010100001) = -351.0    || 21.566122895178978 = 21.0
"0000010101",-- (1010100010) = -350.0    || 21.798248236493887 = 21.0
"0000010110",-- (1010100011) = -349.0    || 22.032817126919305 = 22.0
"0000010110",-- (1010100100) = -348.0    || 22.269854101535188 = 22.0
"0000010110",-- (1010100101) = -347.0    || 22.509383916079937 = 22.0
"0000010110",-- (1010100110) = -346.0    || 22.75143154837111  = 22.0
"0000010110",-- (1010100111) = -345.0    || 22.99602219972207  = 22.0
"0000010111",-- (1010101000) = -344.0    || 23.24318129635416  = 23.0
"0000010111",-- (1010101001) = -343.0    || 23.492934490804053 = 23.0
"0000010111",-- (1010101010) = -342.0    || 23.74530766332579  = 23.0
"0000011000",-- (1010101011) = -341.0    || 24.000326923287048 = 24.0
"0000011000",-- (1010101100) = -340.0    || 24.258018610559425 = 24.0
"0000011000",-- (1010101101) = -339.0    || 24.518409296901893 = 24.0
"0000011000",-- (1010101110) = -338.0    || 24.781525787337397 = 24.0
"0000011001",-- (1010101111) = -337.0    || 25.047395121521767 = 25.0
"0000011001",-- (1010110000) = -336.0    || 25.316044575104634 = 25.0
"0000011001",-- (1010110001) = -335.0    || 25.587501661081934 = 25.0
"0000011001",-- (1010110010) = -334.0    || 25.8617941311392   = 25.0
"0000011010",-- (1010110011) = -333.0    || 26.138949976985504 = 26.0
"0000011010",-- (1010110100) = -332.0    || 26.418997431677234 = 26.0
"0000011010",-- (1010110101) = -331.0    || 26.70196497093117  = 26.0
"0000011010",-- (1010110110) = -330.0    || 26.987881314426637 = 26.0
"0000011011",-- (1010110111) = -329.0    || 27.276775427095664 = 27.0
"0000011011",-- (1010111000) = -328.0    || 27.568676520401027 = 27.0
"0000011011",-- (1010111001) = -327.0    || 27.863614053601285 = 27.0
"0000011100",-- (1010111010) = -326.0    || 28.161617735002338 = 28.0
"0000011100",-- (1010111011) = -325.0    || 28.46271752319495  = 28.0
"0000011100",-- (1010111100) = -324.0    || 28.766943628277357 = 28.0
"0000011101",-- (1010111101) = -323.0    || 29.07432651306266  = 29.0
"0000011101",-- (1010111110) = -322.0    || 29.384896894270103 = 29.0
"0000011101",-- (1010111111) = -321.0    || 29.698685743699578 = 29.0
"0000011110",-- (1011000000) = -320.0    || 30.01572428938887  = 30.0
"0000011110",-- (1011000001) = -319.0    || 30.336044016752723 = 30.0
"0000011110",-- (1011000010) = -318.0    || 30.659676669703053 = 30.0
"0000011110",-- (1011000011) = -317.0    || 30.98665425174983  = 30.0
"0000011111",-- (1011000100) = -316.0    || 31.31700902708143  = 31.0
"0000011111",-- (1011000101) = -315.0    || 31.650773521624238 = 31.0
"0000011111",-- (1011000110) = -314.0    || 31.98798052408026  = 31.0
"0000100000",-- (1011000111) = -313.0    || 32.32866308694225  = 32.0
"0000100000",-- (1011001000) = -312.0    || 32.672854527485505 = 32.0
"0000100001",-- (1011001001) = -311.0    || 33.020588428735394 = 33.0
"0000100001",-- (1011001010) = -310.0    || 33.37189864040995  = 33.0
"0000100001",-- (1011001011) = -309.0    || 33.72681927983662  = 33.0
"0000100010",-- (1011001100) = -308.0    || 34.085384732842144 = 34.0
"0000100010",-- (1011001101) = -307.0    || 34.44762965461516  = 34.0
"0000100010",-- (1011001110) = -306.0    || 34.813588970539975 = 34.0
"0000100011",-- (1011001111) = -305.0    || 35.18329787700124  = 35.0
"0000100011",-- (1011010000) = -304.0    || 35.55679184215815  = 35.0
"0000100011",-- (1011010001) = -303.0    || 35.93410660668743  = 35.0
"0000100100",-- (1011010010) = -302.0    || 36.315278184494225 = 36.0
"0000100100",-- (1011010011) = -301.0    || 36.7003428633896   = 36.0
"0000100101",-- (1011010100) = -300.0    || 37.08933720573413  = 37.0
"0000100101",-- (1011010101) = -299.0    || 37.482298049046165 = 37.0
"0000100101",-- (1011010110) = -298.0    || 37.879262506573845 = 37.0
"0000100110",-- (1011010111) = -297.0    || 38.28026796783013  = 38.0
"0000100110",-- (1011011000) = -296.0    || 38.68535209908924  = 38.0
"0000100111",-- (1011011001) = -295.0    || 39.09455284384402  = 39.0
"0000100111",-- (1011011010) = -294.0    || 39.507908423222624 = 39.0
"0000100111",-- (1011011011) = -293.0    || 39.925457336363735 = 39.0
"0000101000",-- (1011011100) = -292.0    || 40.347238360749174 = 40.0
"0000101000",-- (1011011101) = -291.0    || 40.77329055249249  = 40.0
"0000101001",-- (1011011110) = -290.0    || 41.2036532465828   = 41.0
"0000101001",-- (1011011111) = -289.0    || 41.63836605708225  = 41.0
"0000101010",-- (1011100000) = -288.0    || 42.077468877276175 = 42.0
"0000101010",-- (1011100001) = -287.0    || 42.52100187977483  = 42.0
"0000101010",-- (1011100010) = -286.0    || 42.96900551656503  = 42.0
"0000101011",-- (1011100011) = -285.0    || 43.42152051901103  = 43.0
"0000101011",-- (1011100100) = -284.0    || 43.878587897802895 = 43.0
"0000101100",-- (1011100101) = -283.0    || 44.340248942851225 = 44.0
"0000101100",-- (1011100110) = -282.0    || 44.80654522312722  = 44.0
"0000101101",-- (1011100111) = -281.0    || 45.2775185864462   = 45.0
"0000101101",-- (1011101000) = -280.0    || 45.75321115919381  = 45.0
"0000101110",-- (1011101001) = -279.0    || 46.233665345993174 = 46.0
"0000101110",-- (1011101010) = -278.0    || 46.71892382931171  = 46.0
"0000101111",-- (1011101011) = -277.0    || 47.20902956900649  = 47.0
"0000101111",-- (1011101100) = -276.0    || 47.70402580180614  = 47.0
"0000110000",-- (1011101101) = -275.0    || 48.203956040728634 = 48.0
"0000110000",-- (1011101110) = -274.0    || 48.70886407443282  = 48.0
"0000110001",-- (1011101111) = -273.0    || 49.218793966502574 = 49.0
"0000110001",-- (1011110000) = -272.0    || 49.73379005466228  = 49.0
"0000110010",-- (1011110001) = -271.0    || 50.253896949921575 = 50.0
"0000110010",-- (1011110010) = -270.0    || 50.779159535648496 = 50.0
"0000110011",-- (1011110011) = -269.0    || 51.309622966569094 = 51.0
"0000110011",-- (1011110100) = -268.0    || 51.84533266769187  = 51.0
"0000110100",-- (1011110101) = -267.0    || 52.386334333156164 = 52.0
"0000110100",-- (1011110110) = -266.0    || 52.93267392500187  = 52.0
"0000110101",-- (1011110111) = -265.0    || 53.48439767185995  = 53.0
"0000110110",-- (1011111000) = -264.0    || 54.041552067561334 = 54.0
"0000110110",-- (1011111001) = -263.0    || 54.60418386966298  = 54.0
"0000110111",-- (1011111010) = -262.0    || 55.17234009788949  = 55.0
"0000110111",-- (1011111011) = -261.0    || 55.746068032488246 = 55.0
"0000111000",-- (1011111100) = -260.0    || 56.32541521249704  = 56.0
"0000111000",-- (1011111101) = -259.0    || 56.91042943392188  = 56.0
"0000111001",-- (1011111110) = -258.0    || 57.501158747823446 = 57.0
"0000111010",-- (1011111111) = -257.0    || 58.09765145831112  = 58.0
"0000111010",-- (1100000000) = -256.0    || 58.699956120441605 = 58.0
"0000111011",-- (1100000001) = -255.0    || 59.30812153802183  = 59.0
"0000111011",-- (1100000010) = -254.0    || 59.92219676131329  = 59.0
"0000111100",-- (1100000011) = -253.0    || 60.54223108463647  = 60.0
"0000111101",-- (1100000100) = -252.0    || 61.16827404387403  = 61.0
"0000111101",-- (1100000101) = -251.0    || 61.80037541386994  = 61.0
"0000111110",-- (1100000110) = -250.0    || 62.43858520572397  = 62.0
"0000111111",-- (1100000111) = -249.0    || 63.08295366397874  = 63.0
"0000111111",-- (1100001000) = -248.0    || 63.733531263698126 = 63.0
"0001000000",-- (1100001001) = -247.0    || 64.39036870743512  = 64.0
"0001000001",-- (1100001010) = -246.0    || 65.0535169220869   = 65.0
"0001000001",-- (1100001011) = -245.0    || 65.7230270556362   = 65.0
"0001000010",-- (1100001100) = -244.0    || 66.39895047377593  = 66.0
"0001000011",-- (1100001101) = -243.0    || 67.08133875641624  = 67.0
"0001000011",-- (1100001110) = -242.0    || 67.77024369407191  = 67.0
"0001000100",-- (1100001111) = -241.0    || 68.46571728412758  = 68.0
"0001000101",-- (1100010000) = -240.0    || 69.1678117269802   = 69.0
"0001000101",-- (1100010001) = -239.0    || 69.87657942205566  = 69.0
"0001000110",-- (1100010010) = -238.0    || 70.59207296369833  = 70.0
"0001000111",-- (1100010011) = -237.0    || 71.3143451369319   = 71.0
"0001001000",-- (1100010100) = -236.0    || 72.04344891308892  = 72.0
"0001001000",-- (1100010101) = -235.0    || 72.77943744530795  = 72.0
"0001001001",-- (1100010110) = -234.0    || 73.52236406389606  = 73.0
"0001001010",-- (1100010111) = -233.0    || 74.27228227155477  = 74.0
"0001001011",-- (1100011000) = -232.0    || 75.02924573846818  = 75.0
"0001001011",-- (1100011001) = -231.0    || 75.79330829725056  = 75.0
"0001001100",-- (1100011010) = -230.0    || 76.56452393775244  = 76.0
"0001001101",-- (1100011011) = -229.0    || 77.34294680172287  = 77.0
"0001001110",-- (1100011100) = -228.0    || 78.12863117732613  = 78.0
"0001001110",-- (1100011101) = -227.0    || 78.92163149351134  = 78.0
"0001001111",-- (1100011110) = -226.0    || 79.72200231423282  = 79.0
"0001010000",-- (1100011111) = -225.0    || 80.52979833251989  = 80.0
"0001010001",-- (1100100000) = -224.0    || 81.34507436439388  = 81.0
"0001010010",-- (1100100001) = -223.0    || 82.16788534263083  = 82.0
"0001010010",-- (1100100010) = -222.0    || 82.9982863103685   = 82.0
"0001010011",-- (1100100011) = -221.0    || 83.8363324145552   = 83.0
"0001010100",-- (1100100100) = -220.0    || 84.68207889923978  = 84.0
"0001010101",-- (1100100101) = -219.0    || 85.53558109870012  = 85.0
"0001010110",-- (1100100110) = -218.0    || 86.39689443040918  = 86.0
"0001010111",-- (1100100111) = -217.0    || 87.26607438783692  = 87.0
"0001011000",-- (1100101000) = -216.0    || 88.1431765330861   = 88.0
"0001011001",-- (1100101001) = -215.0    || 89.02825648936108  = 89.0
"0001011001",-- (1100101010) = -214.0    || 89.92136993326743  = 89.0
"0001011010",-- (1100101011) = -213.0    || 90.8225725869412   = 90.0
"0001011011",-- (1100101100) = -212.0    || 91.73192021000683  = 91.0
"0001011100",-- (1100101101) = -211.0    || 92.64946859136116  = 92.0
"0001011101",-- (1100101110) = -210.0    || 93.57527354078347  = 93.0
"0001011110",-- (1100101111) = -209.0    || 94.50939088036938  = 94.0
"0001011111",-- (1100110000) = -208.0    || 95.45187643578737  = 95.0
"0001100000",-- (1100110001) = -207.0    || 96.4027860273574   = 96.0
"0001100001",-- (1100110010) = -206.0    || 97.36217546094927  = 97.0
"0001100010",-- (1100110011) = -205.0    || 98.33010051870083  = 98.0
"0001100011",-- (1100110100) = -204.0    || 99.3066169495539   = 99.0
"0001100100",-- (1100110101) = -203.0    || 100.29178045960732 = 100.0
"0001100101",-- (1100110110) = -202.0    || 101.28564670228664 = 101.0
"0001100110",-- (1100110111) = -201.0    || 102.2882712683281  = 102.0
"0001100111",-- (1100111000) = -200.0    || 103.29970967557787 = 103.0
"0001101000",-- (1100111001) = -199.0    || 104.32001735860425 = 104.0
"0001101001",-- (1100111010) = -198.0    || 105.34924965812252 = 105.0
"0001101010",-- (1100111011) = -197.0    || 106.38746181023262 = 106.0
"0001101011",-- (1100111100) = -196.0    || 107.43470893546747 = 107.0
"0001101100",-- (1100111101) = -195.0    || 108.4910460276529  = 108.0
"0001101101",-- (1100111110) = -194.0    || 109.55652794257776 = 109.0
"0001101110",-- (1100111111) = -193.0    || 110.63120938647411 = 110.0
"0001101111",-- (1101000000) = -192.0    || 111.71514490430769 = 111.0
"0001110000",-- (1101000001) = -191.0    || 112.80838886787724 = 112.0
"0001110001",-- (1101000010) = -190.0    || 113.91099546372408 = 113.0
"0001110011",-- (1101000011) = -189.0    || 115.02301868085063 = 115.0
"0001110100",-- (1101000100) = -188.0    || 116.1445122982483  = 116.0
"0001110101",-- (1101000101) = -187.0    || 117.27552987223544 = 117.0
"0001110110",-- (1101000110) = -186.0    || 118.41612472360471 = 118.0
"0001110111",-- (1101000111) = -185.0    || 119.56634992458054 = 119.0
"0001111000",-- (1101001000) = -184.0    || 120.72625828558762 = 120.0
"0001111001",-- (1101001001) = -183.0    || 121.89590234182975 = 121.0
"0001111011",-- (1101001010) = -182.0    || 123.07533433968132 = 123.0
"0001111100",-- (1101001011) = -181.0    || 124.26460622289028 = 124.0
"0001111101",-- (1101001100) = -180.0    || 125.46376961859504 = 125.0
"0001111110",-- (1101001101) = -179.0    || 126.67287582315541 = 126.0
"0001111111",-- (1101001110) = -178.0    || 127.89197578779911 = 127.0
"0010000001",-- (1101001111) = -177.0    || 129.12112010408433 = 129.0
"0010000010",-- (1101010000) = -176.0    || 130.36035898918064 = 130.0
"0010000011",-- (1101010001) = -175.0    || 131.60974227096895 = 131.0
"0010000100",-- (1101010010) = -174.0    || 132.8693193729624  = 132.0
"0010000110",-- (1101010011) = -173.0    || 134.13913929904973 = 134.0
"0010000111",-- (1101010100) = -172.0    || 135.4192506180632  = 135.0
"0010001000",-- (1101010101) = -171.0    || 136.70970144817252 = 136.0
"0010001010",-- (1101010110) = -170.0    || 138.0105394411078  = 138.0
"0010001011",-- (1101010111) = -169.0    || 139.32181176621236 = 139.0
"0010001100",-- (1101011000) = -168.0    || 140.6435650943296  = 140.0
"0010001101",-- (1101011001) = -167.0    || 141.97584558152448 = 141.0
"0010001111",-- (1101011010) = -166.0    || 143.31869885264385 = 143.0
"0010010000",-- (1101011011) = -165.0    || 144.67216998471764 = 144.0
"0010010010",-- (1101011100) = -164.0    || 146.03630349020418 = 146.0
"0010010011",-- (1101011101) = -163.0    || 147.41114330008253 = 147.0
"0010010100",-- (1101011110) = -162.0    || 148.7967327467953  = 148.0
"0010010110",-- (1101011111) = -161.0    || 150.19311454704538 = 150.0
"0010010111",-- (1101100000) = -160.0    || 151.60033078445002 = 151.0
"0010011001",-- (1101100001) = -159.0    || 153.01842289205618 = 153.0
"0010011010",-- (1101100010) = -158.0    || 154.44743163472103 = 154.0
"0010011011",-- (1101100011) = -157.0    || 155.8873970913614  = 155.0
"0010011101",-- (1101100100) = -156.0    || 157.33835863707716 = 157.0
"0010011110",-- (1101100101) = -155.0    || 158.80035492515182 = 158.0
"0010100000",-- (1101100110) = -154.0    || 160.27342386893628 = 160.0
"0010100001",-- (1101100111) = -153.0    || 161.75760262361905 = 161.0
"0010100011",-- (1101101000) = -152.0    || 163.25292756788915 = 163.0
"0010100100",-- (1101101001) = -151.0    || 164.75943428549604 = 164.0
"0010100110",-- (1101101010) = -150.0    || 166.27715754671192 = 166.0
"0010100111",-- (1101101011) = -149.0    || 167.80613128970228 = 167.0
"0010101001",-- (1101101100) = -148.0    || 169.34638860180974 = 169.0
"0010101010",-- (1101101101) = -147.0    || 170.8979617007574  = 170.0
"0010101100",-- (1101101110) = -146.0    || 172.4608819157776  = 172.0
"0010101110",-- (1101101111) = -145.0    || 174.03517966867213 = 174.0
"0010101111",-- (1101110000) = -144.0    || 175.6208844548105  = 175.0
"0010110001",-- (1101110001) = -143.0    || 177.21802482407222 = 177.0
"0010110010",-- (1101110010) = -142.0    || 178.82662836174046 = 178.0
"0010110100",-- (1101110011) = -141.0    || 180.44672166935388 = 180.0
"0010110110",-- (1101110100) = -140.0    || 182.07833034552277 = 182.0
"0010110111",-- (1101110101) = -139.0    || 183.72147896671837 = 183.0
"0010111001",-- (1101110110) = -138.0    || 185.3761910680409  = 185.0
"0010111011",-- (1101110111) = -137.0    || 187.04248912397574 = 187.0
"0010111100",-- (1101111000) = -136.0    || 188.72039452914387 = 188.0
"0010111110",-- (1101111001) = -135.0    || 190.40992757905582 = 190.0
"0011000000",-- (1101111010) = -134.0    || 192.11110745087635 = 192.0
"0011000001",-- (1101111011) = -133.0    || 193.82395218420854 = 193.0
"0011000011",-- (1101111100) = -132.0    || 195.54847866190565 = 195.0
"0011000101",-- (1101111101) = -131.0    || 197.2847025909197  = 197.0
"0011000111",-- (1101111110) = -130.0    || 199.03263848319455 = 199.0
"0011001000",-- (1101111111) = -129.0    || 200.792299636614   = 200.0
"0011001010",-- (1110000000) = -128.0    || 202.5636981160123  = 202.0
"0011001100",-- (1110000001) = -127.0    || 204.34684473425781 = 204.0
"0011001110",-- (1110000010) = -126.0    || 206.1417490334183  = 206.0
"0011001111",-- (1110000011) = -125.0    || 207.94841926601748 = 207.0
"0011010001",-- (1110000100) = -124.0    || 209.7668623763937  = 209.0
"0011010011",-- (1110000101) = -123.0    || 211.5970839821685  = 211.0
"0011010101",-- (1110000110) = -122.0    || 213.43908835583719 = 213.0
"0011010111",-- (1110000111) = -121.0    || 215.29287840649008 = 215.0
"0011011001",-- (1110001000) = -120.0    || 217.15845566167584 = 217.0
"0011011011",-- (1110001001) = -119.0    || 219.03582024941622 = 219.0
"0011011100",-- (1110001010) = -118.0    || 220.92497088038314 = 220.0
"0011011110",-- (1110001011) = -117.0    || 222.8259048302495  = 222.0
"0011100000",-- (1110001100) = -116.0    || 224.73861792222314 = 224.0
"0011100010",-- (1110001101) = -115.0    || 226.66310450977585 = 226.0
"0011100100",-- (1110001110) = -114.0    || 228.59935745957804 = 228.0
"0011100110",-- (1110001111) = -113.0    || 230.54736813464967 = 230.0
"0011101000",-- (1110010000) = -112.0    || 232.50712637773978 = 232.0
"0011101010",-- (1110010001) = -111.0    || 234.47862049494418 = 234.0
"0011101100",-- (1110010010) = -110.0    || 236.4618372395743  = 236.0
"0011101110",-- (1110010011) = -109.0    || 238.45676179628757 = 238.0
"0011110000",-- (1110010100) = -108.0    || 240.4633777654902  = 240.0
"0011110010",-- (1110010101) = -107.0    || 242.48166714802605 = 242.0
"0011110100",-- (1110010110) = -106.0    || 244.51161033016027 = 244.0
"0011110110",-- (1110010111) = -105.0    || 246.55318606887144 = 246.0
"0011111000",-- (1110011000) = -104.0    || 248.60637147746303 = 248.0
"0011111010",-- (1110011001) = -103.0    || 250.6711420115055  = 250.0
"0011111100",-- (1110011010) = -102.0    || 252.747471455121   = 252.0
"0011111110",-- (1110011011) = -101.0    || 254.8353319076226  = 254.0
"0100000000",-- (1110011100) = -100.0    || 256.934693770519   = 256.0
"0100000011",-- (1110011101) = -99.0     || 259.0455257348971  = 259.0
"0100000101",-- (1110011110) = -98.0     || 261.1677947691931  = 261.0
"0100000111",-- (1110011111) = -97.0     || 263.30146610736455 = 263.0
"0100001001",-- (1110100000) = -96.0     || 265.44650323747436 = 265.0
"0100001011",-- (1110100001) = -95.0     || 267.6028678906986  = 267.0
"0100001101",-- (1110100010) = -94.0     || 269.7705200307691  = 269.0
"0100001111",-- (1110100011) = -93.0     || 271.94941784386225 = 271.0
"0100010010",-- (1110100100) = -92.0     || 274.1395177289456  = 274.0
"0100010100",-- (1110100101) = -91.0     || 276.34077428859285 = 276.0
"0100010110",-- (1110100110) = -90.0     || 278.5531403202791  = 278.0
"0100011000",-- (1110100111) = -89.0     || 280.776566808166   = 280.0
"0100011011",-- (1110101000) = -88.0     || 283.01100291538927 = 283.0
"0100011101",-- (1110101001) = -87.0     || 285.25639597685716 = 285.0
"0100011111",-- (1110101010) = -86.0     || 287.51269149257325 = 287.0
"0100100001",-- (1110101011) = -85.0     || 289.77983312149047 = 289.0
"0100100100",-- (1110101100) = -84.0     || 292.0577626759095  = 292.0
"0100100110",-- (1110101101) = -83.0     || 294.34642011643    = 294.0
"0100101000",-- (1110101110) = -82.0     || 296.64574354746503 = 296.0
"0100101010",-- (1110101111) = -81.0     || 298.9556692133277  = 298.0
"0100101101",-- (1110110000) = -80.0     || 301.2761314949005  = 301.0
"0100101111",-- (1110110001) = -79.0     || 303.60706290689495 = 303.0
"0100110001",-- (1110110010) = -78.0     || 305.9483940957124  = 305.0
"0100110100",-- (1110110011) = -77.0     || 308.30005383791274 = 308.0
"0100110110",-- (1110110100) = -76.0     || 310.6619690393012  = 310.0
"0100111001",-- (1110110101) = -75.0     || 313.03406473463957 = 313.0
"0100111011",-- (1110110110) = -74.0     || 315.4162640879915  = 315.0
"0100111101",-- (1110110111) = -73.0     || 317.8084883937084  = 317.0
"0101000000",-- (1110111000) = -72.0     || 320.21065707806304 = 320.0
"0101000010",-- (1110111001) = -71.0     || 322.6226877015387  = 322.0
"0101000101",-- (1110111010) = -70.0     || 325.04449596178006 = 325.0
"0101000111",-- (1110111011) = -69.0     || 327.47599569721154 = 327.0
"0101001001",-- (1110111100) = -68.0     || 329.91709889132994 = 329.0
"0101001100",-- (1110111101) = -67.0     || 332.3677156776768  = 332.0
"0101001110",-- (1110111110) = -66.0     || 334.82775434549507 = 334.0
"0101010001",-- (1110111111) = -65.0     || 337.29712134607564 = 337.0
"0101010011",-- (1111000000) = -64.0     || 339.7757212997979  = 339.0
"0101010110",-- (1111000001) = -63.0     || 342.2634570038686  = 342.0
"0101011000",-- (1111000010) = -62.0     || 344.76022944076226 = 344.0
"0101011011",-- (1111000011) = -61.0     || 347.2659377873667  = 347.0
"0101011101",-- (1111000100) = -60.0     || 349.7804794248366  = 349.0
"0101100000",-- (1111000101) = -59.0     || 352.3037499491578  = 352.0
"0101100010",-- (1111000110) = -58.0     || 354.8356431824229  = 354.0
"0101100101",-- (1111000111) = -57.0     || 357.37605118482145 = 357.0
"0101100111",-- (1111001000) = -56.0     || 359.9248642673449  = 359.0
"0101101010",-- (1111001001) = -55.0     || 362.48197100520747 = 362.0
"0101101101",-- (1111001010) = -54.0     || 365.0472582519816  = 365.0
"0101101111",-- (1111001011) = -53.0     || 367.6206111544504  = 367.0
"0101110010",-- (1111001100) = -52.0     || 370.20191316817323 = 370.0
"0101110100",-- (1111001101) = -51.0     || 372.7910460737659  = 372.0
"0101110111",-- (1111001110) = -50.0     || 375.3878899938917  = 375.0
"0101111001",-- (1111001111) = -49.0     || 377.99232341096223 = 377.0
"0101111100",-- (1111010000) = -48.0     || 380.60422318554504 = 380.0
"0101111111",-- (1111010001) = -47.0     || 383.2234645754741  = 383.0
"0110000001",-- (1111010010) = -46.0     || 385.8499212556616  = 385.0
"0110000100",-- (1111010011) = -45.0     || 388.4834653386032  = 388.0
"0110000111",-- (1111010100) = -44.0     || 391.1239673955763  = 391.0
"0110001001",-- (1111010101) = -43.0     || 393.7712964785225  = 393.0
"0110001100",-- (1111010110) = -42.0     || 396.4253201426112  = 396.0
"0110001111",-- (1111010111) = -41.0     || 399.085904469476   = 399.0
"0110010001",-- (1111011000) = -40.0     || 401.75291409111895 = 401.0
"0110010100",-- (1111011001) = -39.0     || 404.4262122144746  = 404.0
"0110010111",-- (1111011010) = -38.0     || 407.10566064662584 = 407.0
"0110011001",-- (1111011011) = -37.0     || 409.7911198206643  = 409.0
"0110011100",-- (1111011100) = -36.0     || 412.4824488221857  = 412.0
"0110011111",-- (1111011101) = -35.0     || 415.1795054164116  = 415.0
"0110100001",-- (1111011110) = -34.0     || 417.8821460759275  = 417.0
"0110100100",-- (1111011111) = -33.0     || 420.5902260090275  = 420.0
"0110100111",-- (1111100000) = -32.0     || 423.30359918865406 = 423.0
"0110101010",-- (1111100001) = -31.0     || 426.02211838192335 = 426.0
"0110101100",-- (1111100010) = -30.0     || 428.7456351802232  = 428.0
"0110101111",-- (1111100011) = -29.0     || 431.4740000298716  = 431.0
"0110110010",-- (1111100100) = -28.0     || 434.20706226332493 = 434.0
"0110110100",-- (1111100101) = -27.0     || 436.94467013092094 = 436.0
"0110110111",-- (1111100110) = -26.0     || 439.68667083314466 = 439.0
"0110111010",-- (1111100111) = -25.0     || 442.43291055340217 = 442.0
"0110111101",-- (1111101000) = -24.0     || 445.18323449128974 = 445.0
"0110111111",-- (1111101001) = -23.0     || 447.9374868963422  = 447.0
"0111000010",-- (1111101010) = -22.0     || 450.69551110224614 = 450.0
"0111000101",-- (1111101011) = -21.0     || 453.45714956150226 = 453.0
"0111001000",-- (1111101100) = -20.0     || 456.22224388052246 = 456.0
"0111001010",-- (1111101101) = -19.0     || 458.99063485514307 = 458.0
"0111001101",-- (1111101110) = -18.0     || 461.76216250654016 = 461.0
"0111010000",-- (1111101111) = -17.0     || 464.5366661175293  = 464.0
"0111010011",-- (1111110000) = -16.0     || 467.3139842692313  = 467.0
"0111010110",-- (1111110001) = -15.0     || 470.0939548780887  = 470.0
"0111011000",-- (1111110010) = -14.0     || 472.8764152332146  = 472.0
"0111011011",-- (1111110011) = -13.0     || 475.66120203405393 = 475.0
"0111011110",-- (1111110100) = -12.0     || 478.4481514283418  = 478.0
"0111100001",-- (1111110101) = -11.0     || 481.23709905033854 = 481.0
"0111100100",-- (1111110110) = -10.0     || 484.0278800593233  = 484.0
"0111100110",-- (1111110111) = -9.0      || 486.82032917832566 = 486.0
"0111101001",-- (1111111000) = -8.0      || 489.61428073308    = 489.0
"0111101100",-- (1111111001) = -7.0      || 492.40956869117826 = 492.0
"0111101111",-- (1111111010) = -6.0      || 495.20602670140465 = 495.0
"0111110010",-- (1111111011) = -5.0      || 498.00348813323217 = 498.0
"0111110100",-- (1111111100) = -4.0      || 500.8017861164602  = 500.0
"0111110111",-- (1111111101) = -3.0      || 503.60075358097447 = 503.0
"0111111010",-- (1111111110) = -2.0      || 506.40022329660667 = 506.0
"0111111101",-- (1111111111) = -1.0      || 509.20002791307746 = 509.0

--	2 => "11111111" , --255
--	3 => "11010101" ,
others => "00000000000"
) ;
begin
---------------
data_out <= myrom(to_integer(unsigned(address))) ;
end architecture ;
