
--https://stackoverflow.com/questions/17579716/implementing-rom-in-xilinx-vhdl
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.numeric_std.all;
----------------
ENTITY ROM_fx_6bitaddr_6width is
generic(addr_heigth : integer := 64; -- store 64 elements
				addr_bits  : integer := 6; -- required bits to store 64 elements
				data_width : integer := 6  -- each element has 6-bits
				);
  PORT (
    address : IN STD_LOGIC_VECTOR(addr_bits - 1 DOWNTO 0);
    data_out : OUT STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0)
  );
END ENTITY;
------------------
architecture arch of ROM_fx_6bitaddr_6width is
	type memory is array ( 0 to addr_heigth-1 ) of std_logic_vector(data_width-1 downto 0 ) ;
	constant myrom : memory := (
--"int_f_x",--(address)  =integer_MAC|| f(x)               = int_f_x 
"100000",-- (000000) = 0.0       || 32.0               = 32.0
"100010",-- (000001) = 1.0       || 34.79287598317305  = 34.0
"100101",-- (000010) = 2.0       || 37.54352505070913  = 37.0
"101000",-- (000011) = 3.0       || 40.21223605090344  = 40.0
"101010",-- (000100) = 4.0       || 42.764017418762634 = 42.0
"101101",-- (000101) = 5.0       || 45.17024178156872  = 45.0
"101111",-- (000110) = 6.0       || 47.40959354765785  = 47.0
"110001",-- (000111) = 7.0       || 49.46830460139127  = 49.0
"110011",-- (001000) = 8.0       || 51.33976886774923  = 51.0
"110101",-- (001001) = 9.0       || 53.023694721574344 = 53.0
"110110",-- (001010) = 10.0      || 54.52497932597188  = 54.0
"110111",-- (001011) = 11.0      || 55.85247756317621  = 55.0
"111001",-- (001100) = 12.0      || 57.01780344348077  = 57.0
"111010",-- (001101) = 13.0      || 58.034257722763286 = 58.0
"111010",-- (001110) = 14.0      || 58.91593285222538  = 58.0
"111011",-- (001111) = 15.0      || 59.67701176706374  = 59.0
"111100",-- (010000) = 16.0      || 60.3312527424724   = 60.0
"111100",-- (010001) = 17.0      || 60.891638121583604 = 60.0
"111101",-- (010010) = 18.0      || 61.37015819517024  = 61.0
"111101",-- (010011) = 19.0      || 61.77770050986511  = 61.0
"111110",-- (010100) = 20.0      || 62.12401723191319  = 62.0
"111110",-- (010101) = 21.0      || 62.41774721405596  = 62.0
"111110",-- (010110) = 22.0      || 62.66647395080445  = 62.0
"111110",-- (010111) = 23.0      || 62.87680496353124  = 62.0
"111111",-- (011000) = 24.0      || 63.05446197163052  = 63.0
"111111",-- (011001) = 25.0      || 63.204374345396104 = 63.0
"111111",-- (011010) = 26.0      || 63.330770801157236 = 63.0
"111111",-- (011011) = 27.0      || 63.437266160660805 = 63.0
"111111",-- (011100) = 28.0      || 63.52694135396596  = 63.0
"111111",-- (011101) = 29.0      || 63.602415801058385 = 63.0
"111111",-- (011110) = 30.0      || 63.665911955612266 = 63.0
"111111",-- (011111) = 31.0      || 63.71931221391279  = 63.0
"000000",-- (100000) = -32.0     || 0.2357913535639033 = 0.0
"000000",-- (100001) = -31.0     || 0.2806877860872123 = 0.0
"000000",-- (100010) = -30.0     || 0.3340880443877374 = 0.0
"000000",-- (100011) = -29.0     || 0.39758419894161373 = 0.0
"000000",-- (100100) = -28.0     || 0.4730586460340465 = 0.0
"000000",-- (100101) = -27.0     || 0.5627338393391951 = 0.0
"000000",-- (100110) = -26.0     || 0.6692291988427566 = 0.0
"000000",-- (100111) = -25.0     || 0.7956256546038925 = 0.0
"000000",-- (101000) = -24.0     || 0.9455380283694763 = 0.0
"000001",-- (101001) = -23.0     || 1.1231950364687608 = 1.0
"000001",-- (101010) = -22.0     || 1.3335260491955476 = 1.0
"000001",-- (101011) = -21.0     || 1.5822527859440396 = 1.0
"000001",-- (101100) = -20.0     || 1.8759827680868044 = 1.0
"000010",-- (101101) = -19.0     || 2.2222994901348843 = 2.0
"000010",-- (101110) = -18.0     || 2.629841804829761  = 2.0
"000011",-- (101111) = -17.0     || 3.1083618784163924 = 3.0
"000011",-- (110000) = -16.0     || 3.6687472575276003 = 3.0
"000100",-- (110001) = -15.0     || 4.322988232936263  = 4.0
"000101",-- (110010) = -14.0     || 5.0840671477746175 = 5.0
"000101",-- (110011) = -13.0     || 5.965742277236711  = 5.0
"000110",-- (110100) = -12.0     || 6.982196556519231  = 6.0
"001000",-- (110101) = -11.0     || 8.14752243682379   = 8.0
"001001",-- (110110) = -10.0     || 9.475020674028126  = 9.0
"001010",-- (110111) = -9.0      || 10.976305278425656 = 10.0
"001100",-- (111000) = -8.0      || 12.660231132250768 = 12.0
"001110",-- (111001) = -7.0      || 14.531695398608736 = 14.0
"010000",-- (111010) = -6.0      || 16.590406452342148 = 16.0
"010010",-- (111011) = -5.0      || 18.82975821843128  = 18.0
"010101",-- (111100) = -4.0      || 21.23598258123737  = 21.0
"010111",-- (111101) = -3.0      || 23.787763949096565 = 23.0
"011010",-- (111110) = -2.0      || 26.45647494929088  = 26.0
"011101",-- (111111) = -1.0      || 29.207124016826956 = 29.0

--	2 => "11111111" , --255
--	3 => "11010101" ,
others => "00000000000"
) ;
begin
---------------
data_out <= myrom(to_integer(unsigned(address))) ;
end architecture ;
