

--https://stackoverflow.com/questions/17579716/implementing-rom-in-xilinx-vhdl
LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
use ieee.numeric_std.all;

----------------

ENTITY ROM_fixedpoint_8bit is
generic(addr_width : integer := 256; -- store 256 elements
				addr_bits  : integer := 8; -- required bits to store 256 elements
				data_width : integer := 7  -- each element has 7-bits
				);
			
  PORT (
    address : IN STD_LOGIC_VECTOR(addr_bits - 1 DOWNTO 0);
    data_out : OUT STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0)
  );
END ENTITY;

------------------
architecture arch of ROM_fixedpoint_8bit is

	type memory is array ( 0 to addr_width-1 ) of std_logic_vector(data_width-1 downto 0 ) ;
	constant myrom : memory := (
	
--"bin_data",--(address)MAC     =integer_MAC|| f(x)               = integer_f_x 
"01000000",-- (00000000)0.0        = 0.0    || 0.5                = 64.0
"01000001",-- (00000010)0.0078125  = 2.0    || 0.5124973964842103 = 65.0
"01000011",-- (00000100)0.015625   = 4.0    || 0.52497918747894   = 67.0
"01000100",-- (00000110)0.0234375  = 6.0    || 0.5374298453437496 = 68.0
"01000110",-- (00001000)0.03125    = 8.0    || 0.549833997312478  = 70.0
"01000111",-- (00001010)0.0390625  = 10.0   || 0.5621765008857981 = 71.0
"01001001",-- (00001100)0.046875   = 12.0   || 0.574442516811659  = 73.0
"01001011",-- (00001110)0.0546875  = 14.0   || 0.5866175789173301 = 75.0
"01001100",-- (00010000)0.0625     = 16.0   || 0.598687660112452  = 76.0
"01001110",-- (00010010)0.0703125  = 18.0   || 0.610639233949222  = 78.0
"01001111",-- (00010100)0.078125   = 20.0   || 0.6224593312018546 = 79.0
"01010001",-- (00010110)0.0859375  = 22.0   || 0.6341355910108007 = 81.0
"01010010",-- (00011000)0.09375    = 24.0   || 0.6456563062257954 = 82.0
"01010100",-- (00011010)0.1015625  = 26.0   || 0.6570104626734988 = 84.0
"01010101",-- (00011100)0.109375   = 28.0   || 0.6681877721681662 = 85.0
"01010110",-- (00011110)0.1171875  = 30.0   || 0.679178699175393  = 86.0
"01011000",-- (00100000)0.125      = 32.0   || 0.6899744811276125 = 88.0
"01011001",-- (00100010)0.1328125  = 34.0   || 0.700567142473973  = 89.0
"01011011",-- (00100100)0.140625   = 36.0   || 0.7109495026250039 = 91.0
"01011100",-- (00100110)0.1484375  = 38.0   || 0.7211151780228631 = 92.0
"01011101",-- (00101000)0.15625    = 40.0   || 0.7310585786300049 = 93.0
"01011110",-- (00101010)0.1640625  = 42.0   || 0.740774899182154  = 94.0
"01100000",-- (00101100)0.171875   = 44.0   || 0.7502601055951177 = 96.0
"01100001",-- (00101110)0.1796875  = 46.0   || 0.759510916949111  = 97.0
"01100010",-- (00110000)0.1875     = 48.0   || 0.7685247834990178 = 98.0
"01100011",-- (00110010)0.1953125  = 50.0   || 0.7772998611746911 = 99.0
"01100100",-- (00110100)0.203125   = 52.0   || 0.7858349830425586 = 100.0
"01100101",-- (00110110)0.2109375  = 54.0   || 0.7941296281990528 = 101.0
"01100110",-- (00111000)0.21875    = 56.0   || 0.8021838885585818 = 102.0
"01100111",-- (00111010)0.2265625  = 58.0   || 0.8099984339846871 = 103.0
"01101000",-- (00111100)0.234375   = 60.0   || 0.8175744761936437 = 104.0
"01101001",-- (00111110)0.2421875  = 62.0   || 0.8249137318359602 = 105.0
"01101010",-- (01000000)0.25       = 64.0   || 0.8320183851339245 = 106.0
"01101011",-- (01000010)0.2578125  = 66.0   || 0.8388910504234147 = 107.0
"01101100",-- (01000100)0.265625   = 68.0   || 0.8455347349164652 = 108.0
"01101101",-- (01000110)0.2734375  = 70.0   || 0.8519528019683106 = 109.0
"01101101",-- (01001000)0.28125    = 72.0   || 0.8581489350995123 = 109.0
"01101110",-- (01001010)0.2890625  = 74.0   || 0.8641271029909058 = 110.0
"01101111",-- (01001100)0.296875   = 76.0   || 0.8698915256370021 = 111.0
"01110000",-- (01001110)0.3046875  = 78.0   || 0.8754466418125836 = 112.0
"01110000",-- (01010000)0.3125     = 80.0   || 0.8807970779778823 = 112.0
"01110001",-- (01010010)0.3203125  = 82.0   || 0.8859476187202091 = 113.0
"01110010",-- (01010100)0.328125   = 84.0   || 0.8909031788043871 = 114.0
"01110010",-- (01010110)0.3359375  = 86.0   || 0.8956687768809987 = 114.0
"01110011",-- (01011000)0.34375    = 88.0   || 0.9002495108803148 = 115.0
"01110011",-- (01011010)0.3515625  = 90.0   || 0.9046505351008906 = 115.0
"01110100",-- (01011100)0.359375   = 92.0   || 0.9088770389851438 = 116.0
"01110100",-- (01011110)0.3671875  = 94.0   || 0.9129342275597286 = 116.0
"01110101",-- (01100000)0.375      = 96.0   || 0.9168273035060777 = 117.0
"01110101",-- (01100010)0.3828125  = 98.0   || 0.9205614508160216 = 117.0
"01110110",-- (01100100)0.390625   = 100.0  || 0.9241418199787566 = 118.0
"01110110",-- (01100110)0.3984375  = 102.0  || 0.9275735146384823 = 118.0
"01110111",-- (01101000)0.40625    = 104.0  || 0.9308615796566533 = 119.0
"01110111",-- (01101010)0.4140625  = 106.0  || 0.9340109905087812 = 119.0
"01110111",-- (01101100)0.421875   = 108.0  || 0.9370266439430035 = 119.0
"01111000",-- (01101110)0.4296875  = 110.0  || 0.9399133498259924 = 120.0
"01111000",-- (01110000)0.4375     = 112.0  || 0.9426758241011313 = 120.0
"01111001",-- (01110010)0.4453125  = 114.0  || 0.9453186827840592 = 121.0
"01111001",-- (01110100)0.453125   = 116.0  || 0.9478464369215823 = 121.0
"01111001",-- (01110110)0.4609375  = 118.0  || 0.9502634884414434 = 121.0
"01111001",-- (01111000)0.46875    = 120.0  || 0.9525741268224334 = 121.0
"01111010",-- (01111010)0.4765625  = 122.0  || 0.9547825265167125 = 122.0
"01111010",-- (01111100)0.484375   = 124.0  || 0.9568927450589139 = 122.0
"01111010",-- (01111110)0.4921875  = 126.0  || 0.958908721799535  = 122.0
"01111010",-- (01111111)0.5        = 127.0  || 0.9608342772032357 = 122.0
"01111011",-- (01111111)0.5078125  = 127.0  || 0.9626731126558706 = 123.0
"01111011",-- (01111111)0.515625   = 127.0  || 0.9644288107273639 = 123.0
"01111011",-- (01111111)0.5234375  = 127.0  || 0.9661048358408219 = 123.0
"01111011",-- (01111111)0.53125    = 127.0  || 0.9677045353015495 = 123.0
"01111100",-- (01111111)0.5390625  = 127.0  || 0.969231140642852  = 124.0
"01111100",-- (01111111)0.546875   = 127.0  || 0.9706877692486436 = 124.0
"01111100",-- (01111111)0.5546875  = 127.0  || 0.9720774262159271 = 124.0
"01111100",-- (01111111)0.5625     = 127.0  || 0.973403006423134  = 124.0
"01111100",-- (01111111)0.5703125  = 127.0  || 0.9746672967731284 = 124.0
"01111100",-- (01111111)0.578125   = 127.0  || 0.9758729785823308 = 124.0
"01111101",-- (01111111)0.5859375  = 127.0  || 0.9770226300899744 = 125.0
"01111101",-- (01111111)0.59375    = 127.0  || 0.9781187290638694 = 125.0
"01111101",-- (01111111)0.6015625  = 127.0  || 0.9791636554813196 = 125.0
"01111101",-- (01111111)0.609375   = 127.0  || 0.9801596942659225 = 125.0
"01111101",-- (01111111)0.6171875  = 127.0  || 0.9811090380629609 = 125.0
"01111101",-- (01111111)0.625      = 127.0  || 0.9820137900379085 = 125.0
"01111101",-- (01111111)0.6328125  = 127.0  || 0.9828759666842724 = 125.0
"01111101",-- (01111111)0.640625   = 127.0  || 0.9836975006285591 = 125.0
"01111110",-- (01111111)0.6484375  = 127.0  || 0.9844802434215911 = 126.0
"01111110",-- (01111111)0.65625    = 127.0  || 0.9852259683067269 = 126.0
"01111110",-- (01111111)0.6640625  = 127.0  || 0.9859363729567544 = 126.0
"01111110",-- (01111111)0.671875   = 127.0  || 0.9866130821723351 = 126.0
"01111110",-- (01111111)0.6796875  = 127.0  || 0.9872576505358884 = 126.0
"01111110",-- (01111111)0.6875     = 127.0  || 0.9878715650157257 = 126.0
"01111110",-- (01111111)0.6953125  = 127.0  || 0.9884562475160777 = 126.0
"01111110",-- (01111111)0.703125   = 127.0  || 0.9890130573694068 = 126.0
"01111110",-- (01111111)0.7109375  = 127.0  || 0.9895432937680818 = 126.0
"01111110",-- (01111111)0.71875    = 127.0  || 0.9900481981330957 = 126.0
"01111110",-- (01111111)0.7265625  = 127.0  || 0.9905289564180538 = 126.0
"01111110",-- (01111111)0.734375   = 127.0  || 0.990986701347152  = 126.0
"01111110",-- (01111111)0.7421875  = 127.0  || 0.991422514586288  = 126.0
"01111110",-- (01111111)0.75       = 127.0  || 0.9918374288468401 = 126.0
"01111111",-- (01111111)0.7578125  = 127.0  || 0.9922324299219849 = 127.0
"01111111",-- (01111111)0.765625   = 127.0  || 0.9926084586557181 = 127.0
"01111111",-- (01111111)0.7734375  = 127.0  || 0.9929664128450049 = 127.0
"01111111",-- (01111111)0.78125    = 127.0  || 0.9933071490757153 = 127.0
"01111111",-- (01111111)0.7890625  = 127.0  || 0.9936314844931846 = 127.0
"01111111",-- (01111111)0.796875   = 127.0  || 0.9939401985084158 = 127.0
"01111111",-- (01111111)0.8046875  = 127.0  || 0.994234034441075  = 127.0
"01111111",-- (01111111)0.8125     = 127.0  || 0.9945137011005495 = 127.0
"01111111",-- (01111111)0.8203125  = 127.0  || 0.9947798743064417 = 127.0
"01111111",-- (01111111)0.828125   = 127.0  || 0.995033198349943  = 127.0
"01111111",-- (01111111)0.8359375  = 127.0  || 0.9952742873976046 = 127.0
"01111111",-- (01111111)0.84375    = 127.0  || 0.9955037268390589 = 127.0
"01111111",-- (01111111)0.8515625  = 127.0  || 0.9957220745802952 = 127.0
"01111111",-- (01111111)0.859375   = 127.0  || 0.995929862284104  = 127.0
"01111111",-- (01111111)0.8671875  = 127.0  || 0.9961275965593289 = 127.0
"01111111",-- (01111111)0.875      = 127.0  || 0.9963157601005641 = 127.0
"01111111",-- (01111111)0.8828125  = 127.0  || 0.9964948127799336 = 127.0
"01111111",-- (01111111)0.890625   = 127.0  || 0.9966651926925867 = 127.0
"01111111",-- (01111111)0.8984375  = 127.0  || 0.9968273171575148 = 127.0
"01111111",-- (01111111)0.90625    = 127.0  || 0.9969815836752917 = 127.0
"01111111",-- (01111111)0.9140625  = 127.0  || 0.9971283708442995 = 127.0
"01111111",-- (01111111)0.921875   = 127.0  || 0.997268039236989  = 127.0
"01111111",-- (01111111)0.9296875  = 127.0  || 0.9974009322376768 = 127.0
"01111111",-- (01111111)0.9375     = 127.0  || 0.9975273768433653 = 127.0
"01111111",-- (01111111)0.9453125  = 127.0  || 0.997647684429022  = 127.0
"01111111",-- (01111111)0.953125   = 127.0  || 0.9977621514787236 = 127.0
"01111111",-- (01111111)0.9609375  = 127.0  || 0.9978710602840357 = 127.0
"01111111",-- (01111111)0.96875    = 127.0  || 0.9979746796109501 = 127.0
"01111111",-- (01111111)0.9765625  = 127.0  || 0.9980732653366725 = 127.0
"01111111",-- (01111111)0.984375   = 127.0  || 0.9981670610575072 = 127.0
"01111111",-- (01111111)0.9921875  = 127.0  || 0.9982562986690452 = 127.0
"00000000",-- (10000000)-1.0       = -128.0 || 0.0016588010801744215 = 0.0
"00000000",-- (10000000)-0.9921875 = -128.0 || 0.001743701330954778 = 0.0
"00000000",-- (10000000)-0.984375  = -128.0 || 0.0018329389424928035 = 0.0
"00000000",-- (10000000)-0.9765625 = -128.0 || 0.0019267346633274757 = 0.0
"00000000",-- (10000000)-0.96875   = -128.0 || 0.002025320389049882 = 0.0
"00000000",-- (10000000)-0.9609375 = -128.0 || 0.0021289397159641892 = 0.0
"00000000",-- (10000000)-0.953125  = -128.0 || 0.0022378485212763317 = 0.0
"00000000",-- (10000000)-0.9453125 = -128.0 || 0.0023523155709781456 = 0.0
"00000000",-- (10000000)-0.9375    = -128.0 || 0.0024726231566347743 = 0.0
"00000000",-- (10000000)-0.9296875 = -128.0 || 0.002599067762323347 = 0.0
"00000000",-- (10000000)-0.921875  = -128.0 || 0.002731960763011059 = 0.0
"00000000",-- (10000000)-0.9140625 = -128.0 || 0.0028716291557003976 = 0.0
"00000000",-- (10000000)-0.90625   = -128.0 || 0.0030184163247084215 = 0.0
"00000000",-- (10000000)-0.8984375 = -128.0 || 0.0031726828424851893 = 0.0
"00000000",-- (10000000)-0.890625  = -128.0 || 0.0033348073074133443 = 0.0
"00000000",-- (10000000)-0.8828125 = -128.0 || 0.003505187220066338 = 0.0
"00000000",-- (10000000)-0.875     = -128.0 || 0.003684239899435986 = 0.0
"00000000",-- (10000000)-0.8671875 = -128.0 || 0.0038724034406710283 = 0.0
"00000000",-- (10000000)-0.859375  = -128.0 || 0.004070137715896128 = 0.0
"00000000",-- (10000000)-0.8515625 = -128.0 || 0.004277925419704973 = 0.0
"00000000",-- (10000000)-0.84375   = -128.0 || 0.004496273160941178 = 0.0
"00000000",-- (10000000)-0.8359375 = -128.0 || 0.004725712602395478 = 0.0
"00000000",-- (10000000)-0.828125  = -128.0 || 0.004966801650056957 = 0.0
"00000000",-- (10000000)-0.8203125 = -128.0 || 0.005220125693558397 = 0.0
"00000000",-- (10000000)-0.8125    = -128.0 || 0.005486298899450404 = 0.0
"00000000",-- (10000000)-0.8046875 = -128.0 || 0.005765965558924903 = 0.0
"00000000",-- (10000000)-0.796875  = -128.0 || 0.00605980149158411 = 0.0
"00000000",-- (10000000)-0.7890625 = -128.0 || 0.006368515506815542 = 0.0
"00000000",-- (10000000)-0.78125   = -128.0 || 0.0066928509242848554 = 0.0
"00000000",-- (10000000)-0.7734375 = -128.0 || 0.007033587154995161 = 0.0
"00000000",-- (10000000)-0.765625  = -128.0 || 0.007391541344281971 = 0.0
"00000000",-- (10000000)-0.7578125 = -128.0 || 0.007767570078014998 = 0.0
"00000001",-- (10000000)-0.75      = -128.0 || 0.00816257115315989 = 1.0
"00000001",-- (10000000)-0.7421875 = -128.0 || 0.008577485413711984 = 1.0
"00000001",-- (10000000)-0.734375  = -128.0 || 0.009013298652847822 = 1.0
"00000001",-- (10000000)-0.7265625 = -128.0 || 0.009471043581946108 = 1.0
"00000001",-- (10000000)-0.71875   = -128.0 || 0.009951801866904317 = 1.0
"00000001",-- (10000000)-0.7109375 = -128.0 || 0.010456706231918071 = 1.0
"00000001",-- (10000000)-0.703125  = -128.0 || 0.01098694263059318 = 1.0
"00000001",-- (10000000)-0.6953125 = -128.0 || 0.011543752483922289 = 1.0
"00000001",-- (10000000)-0.6875    = -128.0 || 0.012128434984274237 = 1.0
"00000001",-- (10000000)-0.6796875 = -128.0 || 0.012742349464111596 = 1.0
"00000001",-- (10000000)-0.671875  = -128.0 || 0.013386917827664779 = 1.0
"00000001",-- (10000000)-0.6640625 = -128.0 || 0.014063627043245475 = 1.0
"00000001",-- (10000000)-0.65625   = -128.0 || 0.014774031693273055 = 1.0
"00000001",-- (10000000)-0.6484375 = -128.0 || 0.015519756578408886 = 1.0
"00000010",-- (10000000)-0.640625  = -128.0 || 0.01630249937144093 = 2.0
"00000010",-- (10000000)-0.6328125 = -128.0 || 0.017124033315727736 = 2.0
"00000010",-- (10000000)-0.625     = -128.0 || 0.01798620996209156 = 2.0
"00000010",-- (10000000)-0.6171875 = -128.0 || 0.01889096193703905 = 2.0
"00000010",-- (10000000)-0.609375  = -128.0 || 0.019840305734077503 = 2.0
"00000010",-- (10000000)-0.6015625 = -128.0 || 0.020836344518680425 = 2.0
"00000010",-- (10000000)-0.59375   = -128.0 || 0.021881270936130466 = 2.0
"00000010",-- (10000000)-0.5859375 = -128.0 || 0.022977369910025615 = 2.0
"00000011",-- (10000000)-0.578125  = -128.0 || 0.024127021417669196 = 3.0
"00000011",-- (10000000)-0.5703125 = -128.0 || 0.02533270322687172 = 3.0
"00000011",-- (10000000)-0.5625    = -128.0 || 0.026596993576865856 = 3.0
"00000011",-- (10000000)-0.5546875 = -128.0 || 0.027922573784073014 = 3.0
"00000011",-- (10000000)-0.546875  = -128.0 || 0.02931223075135632 = 3.0
"00000011",-- (10000000)-0.5390625 = -128.0 || 0.030768859357148008 = 3.0
"00000100",-- (10000000)-0.53125   = -128.0 || 0.032295464698450495 = 4.0
"00000100",-- (10000000)-0.5234375 = -128.0 || 0.03389516415917814 = 4.0
"00000100",-- (10000000)-0.515625  = -128.0 || 0.03557118927263617 = 4.0
"00000100",-- (10000000)-0.5078125 = -128.0 || 0.03732688734412946 = 4.0
"00000101",-- (10000000)-0.5       = -128.0 || 0.039165722796764356 = 5.0
"00000101",-- (10000010)-0.4921875 = -126.0 || 0.041091278200464994 = 5.0
"00000101",-- (10000100)-0.484375  = -124.0 || 0.043107254941086116 = 5.0
"00000101",-- (10000110)-0.4765625 = -122.0 || 0.04521747348328748 = 5.0
"00000110",-- (10001000)-0.46875   = -120.0 || 0.04742587317756678 = 6.0
"00000110",-- (10001010)-0.4609375 = -118.0 || 0.04973651155855672 = 6.0
"00000110",-- (10001100)-0.453125  = -116.0 || 0.05215356307841772 = 6.0
"00000110",-- (10001110)-0.4453125 = -114.0 || 0.05468131721594076 = 6.0
"00000111",-- (10010000)-0.4375    = -112.0 || 0.05732417589886873 = 7.0
"00000111",-- (10010010)-0.4296875 = -110.0 || 0.060086650174007626 = 7.0
"00001000",-- (10010100)-0.421875  = -108.0 || 0.06297335605699649 = 8.0
"00001000",-- (10010110)-0.4140625 = -106.0 || 0.06598900949121876 = 8.0
"00001000",-- (10011000)-0.40625   = -104.0 || 0.06913842034334682 = 8.0
"00001001",-- (10011010)-0.3984375 = -102.0 || 0.07242648536151769 = 9.0
"00001001",-- (10011100)-0.390625  = -100.0 || 0.07585818002124355 = 9.0
"00001010",-- (10011110)-0.3828125 = -98.0  || 0.07943854918397836 = 10.0
"00001010",-- (10100000)-0.375     = -96.0  || 0.08317269649392235 = 10.0
"00001011",-- (10100010)-0.3671875 = -94.0  || 0.08706577244027125 = 11.0
"00001011",-- (10100100)-0.359375  = -92.0  || 0.09112296101485612 = 11.0
"00001100",-- (10100110)-0.3515625 = -90.0  || 0.09534946489910949 = 12.0
"00001100",-- (10101000)-0.34375   = -88.0  || 0.09975048911968513 = 12.0
"00001101",-- (10101010)-0.3359375 = -86.0  || 0.10433122311900131 = 13.0
"00001101",-- (10101100)-0.328125  = -84.0  || 0.10909682119561294 = 13.0
"00001110",-- (10101110)-0.3203125 = -82.0  || 0.11405238127979084 = 14.0
"00001111",-- (10110000)-0.3125    = -80.0  || 0.11920292202211755 = 15.0
"00001111",-- (10110010)-0.3046875 = -78.0  || 0.12455335818741639 = 15.0
"00010000",-- (10110100)-0.296875  = -76.0  || 0.13010847436299783 = 16.0
"00010001",-- (10110110)-0.2890625 = -74.0  || 0.13587289700909427 = 17.0
"00010010",-- (10111000)-0.28125   = -72.0  || 0.14185106490048777 = 18.0
"00010010",-- (10111010)-0.2734375 = -70.0  || 0.14804719803168948 = 18.0
"00010011",-- (10111100)-0.265625  = -68.0  || 0.15446526508353467 = 19.0
"00010100",-- (10111110)-0.2578125 = -66.0  || 0.16110894957658523 = 20.0
"00010101",-- (11000000)-0.25      = -64.0  || 0.16798161486607552 = 21.0
"00010110",-- (11000010)-0.2421875 = -62.0  || 0.1750862681640398 = 22.0
"00010111",-- (11000100)-0.234375  = -60.0  || 0.18242552380635635 = 23.0
"00011000",-- (11000110)-0.2265625 = -58.0  || 0.19000156601531293 = 24.0
"00011001",-- (11001000)-0.21875   = -56.0  || 0.19781611144141822 = 25.0
"00011010",-- (11001010)-0.2109375 = -54.0  || 0.20587037180094733 = 26.0
"00011011",-- (11001100)-0.203125  = -52.0  || 0.2141650169574414 = 27.0
"00011100",-- (11001110)-0.1953125 = -50.0  || 0.22270013882530884 = 28.0
"00011101",-- (11010000)-0.1875    = -48.0  || 0.23147521650098232 = 29.0
"00011110",-- (11010010)-0.1796875 = -46.0  || 0.24048908305088887 = 30.0
"00011111",-- (11010100)-0.171875  = -44.0  || 0.24973989440488234 = 31.0
"00100001",-- (11010110)-0.1640625 = -42.0  || 0.259225100817846  = 33.0
"00100010",-- (11011000)-0.15625   = -40.0  || 0.2689414213699951 = 34.0
"00100011",-- (11011010)-0.1484375 = -38.0  || 0.2788848219771369 = 35.0
"00100100",-- (11011100)-0.140625  = -36.0  || 0.289050497374996  = 36.0
"00100110",-- (11011110)-0.1328125 = -34.0  || 0.29943285752602705 = 38.0
"00100111",-- (11100000)-0.125     = -32.0  || 0.31002551887238755 = 39.0
"00101001",-- (11100010)-0.1171875 = -30.0  || 0.320821300824607  = 41.0
"00101010",-- (11100100)-0.109375  = -28.0  || 0.3318122278318339 = 42.0
"00101011",-- (11100110)-0.1015625 = -26.0  || 0.34298953732650117 = 43.0
"00101101",-- (11101000)-0.09375   = -24.0  || 0.35434369377420455 = 45.0
"00101110",-- (11101010)-0.0859375 = -22.0  || 0.36586440898919936 = 46.0
"00110000",-- (11101100)-0.078125  = -20.0  || 0.3775406687981454 = 48.0
"00110001",-- (11101110)-0.0703125 = -18.0  || 0.389360766050778  = 49.0
"00110011",-- (11110000)-0.0625    = -16.0  || 0.401312339887548  = 51.0
"00110100",-- (11110010)-0.0546875 = -14.0  || 0.41338242108267   = 52.0
"00110110",-- (11110100)-0.046875  = -12.0  || 0.425557483188341  = 54.0
"00111000",-- (11110110)-0.0390625 = -10.0  || 0.43782349911420193 = 56.0
"00111001",-- (11111000)-0.03125   = -8.0   || 0.45016600268752216 = 57.0
"00111011",-- (11111010)-0.0234375 = -6.0   || 0.46257015465625045 = 59.0
"00111100",-- (11111100)-0.015625  = -4.0   || 0.47502081252106   = 60.0
"00111110",-- (11111110)-0.0078125 = -2.0   || 0.4875026035157896 = 62.0

	
--	2 => "11111111" , --255
--	3 => "11010101" ,  
others => "00000000000" 
) ;

begin 
---------------
data_out <= myrom(to_integer(unsigned(address))) ;
end architecture ;

