LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada2_ReLU_30neuron_8bits_50n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c2_n0_bias, c2_n1_bias, c2_n2_bias, c2_n3_bias, c2_n4_bias, c2_n5_bias, c2_n6_bias, c2_n7_bias, c2_n8_bias, c2_n9_bias, c2_n10_bias, c2_n11_bias, c2_n12_bias, c2_n13_bias, c2_n14_bias, c2_n15_bias, c2_n16_bias, c2_n17_bias, c2_n18_bias, c2_n19_bias, c2_n20_bias, c2_n21_bias, c2_n22_bias, c2_n23_bias, c2_n24_bias, c2_n25_bias, c2_n26_bias, c2_n27_bias, c2_n28_bias, c2_n29_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, c2_n0_w1, c2_n0_w2, c2_n0_w3, c2_n0_w4, c2_n0_w5, c2_n0_w6, c2_n0_w7, c2_n0_w8, c2_n0_w9, c2_n0_w10, c2_n0_w11, c2_n0_w12, c2_n0_w13, c2_n0_w14, c2_n0_w15, c2_n0_w16, c2_n0_w17, c2_n0_w18, c2_n0_w19, c2_n0_w20, c2_n0_w21, c2_n0_w22, c2_n0_w23, c2_n0_w24, c2_n0_w25, c2_n0_w26, c2_n0_w27, c2_n0_w28, c2_n0_w29, c2_n0_w30, c2_n0_w31, c2_n0_w32, c2_n0_w33, c2_n0_w34, c2_n0_w35, c2_n0_w36, c2_n0_w37, c2_n0_w38, c2_n0_w39, c2_n0_w40, c2_n0_w41, c2_n0_w42, c2_n0_w43, c2_n0_w44, c2_n0_w45, c2_n0_w46, c2_n0_w47, c2_n0_w48, c2_n0_w49, c2_n0_w50, c2_n1_w1, c2_n1_w2, c2_n1_w3, c2_n1_w4, c2_n1_w5, c2_n1_w6, c2_n1_w7, c2_n1_w8, c2_n1_w9, c2_n1_w10, c2_n1_w11, c2_n1_w12, c2_n1_w13, c2_n1_w14, c2_n1_w15, c2_n1_w16, c2_n1_w17, c2_n1_w18, c2_n1_w19, c2_n1_w20, c2_n1_w21, c2_n1_w22, c2_n1_w23, c2_n1_w24, c2_n1_w25, c2_n1_w26, c2_n1_w27, c2_n1_w28, c2_n1_w29, c2_n1_w30, c2_n1_w31, c2_n1_w32, c2_n1_w33, c2_n1_w34, c2_n1_w35, c2_n1_w36, c2_n1_w37, c2_n1_w38, c2_n1_w39, c2_n1_w40, c2_n1_w41, c2_n1_w42, c2_n1_w43, c2_n1_w44, c2_n1_w45, c2_n1_w46, c2_n1_w47, c2_n1_w48, c2_n1_w49, c2_n1_w50, c2_n2_w1, c2_n2_w2, c2_n2_w3, c2_n2_w4, c2_n2_w5, c2_n2_w6, c2_n2_w7, c2_n2_w8, c2_n2_w9, c2_n2_w10, c2_n2_w11, c2_n2_w12, c2_n2_w13, c2_n2_w14, c2_n2_w15, c2_n2_w16, c2_n2_w17, c2_n2_w18, c2_n2_w19, c2_n2_w20, c2_n2_w21, c2_n2_w22, c2_n2_w23, c2_n2_w24, c2_n2_w25, c2_n2_w26, c2_n2_w27, c2_n2_w28, c2_n2_w29, c2_n2_w30, c2_n2_w31, c2_n2_w32, c2_n2_w33, c2_n2_w34, c2_n2_w35, c2_n2_w36, c2_n2_w37, c2_n2_w38, c2_n2_w39, c2_n2_w40, c2_n2_w41, c2_n2_w42, c2_n2_w43, c2_n2_w44, c2_n2_w45, c2_n2_w46, c2_n2_w47, c2_n2_w48, c2_n2_w49, c2_n2_w50, c2_n3_w1, c2_n3_w2, c2_n3_w3, c2_n3_w4, c2_n3_w5, c2_n3_w6, c2_n3_w7, c2_n3_w8, c2_n3_w9, c2_n3_w10, c2_n3_w11, c2_n3_w12, c2_n3_w13, c2_n3_w14, c2_n3_w15, c2_n3_w16, c2_n3_w17, c2_n3_w18, c2_n3_w19, c2_n3_w20, c2_n3_w21, c2_n3_w22, c2_n3_w23, c2_n3_w24, c2_n3_w25, c2_n3_w26, c2_n3_w27, c2_n3_w28, c2_n3_w29, c2_n3_w30, c2_n3_w31, c2_n3_w32, c2_n3_w33, c2_n3_w34, c2_n3_w35, c2_n3_w36, c2_n3_w37, c2_n3_w38, c2_n3_w39, c2_n3_w40, c2_n3_w41, c2_n3_w42, c2_n3_w43, c2_n3_w44, c2_n3_w45, c2_n3_w46, c2_n3_w47, c2_n3_w48, c2_n3_w49, c2_n3_w50, c2_n4_w1, c2_n4_w2, c2_n4_w3, c2_n4_w4, c2_n4_w5, c2_n4_w6, c2_n4_w7, c2_n4_w8, c2_n4_w9, c2_n4_w10, c2_n4_w11, c2_n4_w12, c2_n4_w13, c2_n4_w14, c2_n4_w15, c2_n4_w16, c2_n4_w17, c2_n4_w18, c2_n4_w19, c2_n4_w20, c2_n4_w21, c2_n4_w22, c2_n4_w23, c2_n4_w24, c2_n4_w25, c2_n4_w26, c2_n4_w27, c2_n4_w28, c2_n4_w29, c2_n4_w30, c2_n4_w31, c2_n4_w32, c2_n4_w33, c2_n4_w34, c2_n4_w35, c2_n4_w36, c2_n4_w37, c2_n4_w38, c2_n4_w39, c2_n4_w40, c2_n4_w41, c2_n4_w42, c2_n4_w43, c2_n4_w44, c2_n4_w45, c2_n4_w46, c2_n4_w47, c2_n4_w48, c2_n4_w49, c2_n4_w50, c2_n5_w1, c2_n5_w2, c2_n5_w3, c2_n5_w4, c2_n5_w5, c2_n5_w6, c2_n5_w7, c2_n5_w8, c2_n5_w9, c2_n5_w10, c2_n5_w11, c2_n5_w12, c2_n5_w13, c2_n5_w14, c2_n5_w15, c2_n5_w16, c2_n5_w17, c2_n5_w18, c2_n5_w19, c2_n5_w20, c2_n5_w21, c2_n5_w22, c2_n5_w23, c2_n5_w24, c2_n5_w25, c2_n5_w26, c2_n5_w27, c2_n5_w28, c2_n5_w29, c2_n5_w30, c2_n5_w31, c2_n5_w32, c2_n5_w33, c2_n5_w34, c2_n5_w35, c2_n5_w36, c2_n5_w37, c2_n5_w38, c2_n5_w39, c2_n5_w40, c2_n5_w41, c2_n5_w42, c2_n5_w43, c2_n5_w44, c2_n5_w45, c2_n5_w46, c2_n5_w47, c2_n5_w48, c2_n5_w49, c2_n5_w50, c2_n6_w1, c2_n6_w2, c2_n6_w3, c2_n6_w4, c2_n6_w5, c2_n6_w6, c2_n6_w7, c2_n6_w8, c2_n6_w9, c2_n6_w10, c2_n6_w11, c2_n6_w12, c2_n6_w13, c2_n6_w14, c2_n6_w15, c2_n6_w16, c2_n6_w17, c2_n6_w18, c2_n6_w19, c2_n6_w20, c2_n6_w21, c2_n6_w22, c2_n6_w23, c2_n6_w24, c2_n6_w25, c2_n6_w26, c2_n6_w27, c2_n6_w28, c2_n6_w29, c2_n6_w30, c2_n6_w31, c2_n6_w32, c2_n6_w33, c2_n6_w34, c2_n6_w35, c2_n6_w36, c2_n6_w37, c2_n6_w38, c2_n6_w39, c2_n6_w40, c2_n6_w41, c2_n6_w42, c2_n6_w43, c2_n6_w44, c2_n6_w45, c2_n6_w46, c2_n6_w47, c2_n6_w48, c2_n6_w49, c2_n6_w50, c2_n7_w1, c2_n7_w2, c2_n7_w3, c2_n7_w4, c2_n7_w5, c2_n7_w6, c2_n7_w7, c2_n7_w8, c2_n7_w9, c2_n7_w10, c2_n7_w11, c2_n7_w12, c2_n7_w13, c2_n7_w14, c2_n7_w15, c2_n7_w16, c2_n7_w17, c2_n7_w18, c2_n7_w19, c2_n7_w20, c2_n7_w21, c2_n7_w22, c2_n7_w23, c2_n7_w24, c2_n7_w25, c2_n7_w26, c2_n7_w27, c2_n7_w28, c2_n7_w29, c2_n7_w30, c2_n7_w31, c2_n7_w32, c2_n7_w33, c2_n7_w34, c2_n7_w35, c2_n7_w36, c2_n7_w37, c2_n7_w38, c2_n7_w39, c2_n7_w40, c2_n7_w41, c2_n7_w42, c2_n7_w43, c2_n7_w44, c2_n7_w45, c2_n7_w46, c2_n7_w47, c2_n7_w48, c2_n7_w49, c2_n7_w50, c2_n8_w1, c2_n8_w2, c2_n8_w3, c2_n8_w4, c2_n8_w5, c2_n8_w6, c2_n8_w7, c2_n8_w8, c2_n8_w9, c2_n8_w10, c2_n8_w11, c2_n8_w12, c2_n8_w13, c2_n8_w14, c2_n8_w15, c2_n8_w16, c2_n8_w17, c2_n8_w18, c2_n8_w19, c2_n8_w20, c2_n8_w21, c2_n8_w22, c2_n8_w23, c2_n8_w24, c2_n8_w25, c2_n8_w26, c2_n8_w27, c2_n8_w28, c2_n8_w29, c2_n8_w30, c2_n8_w31, c2_n8_w32, c2_n8_w33, c2_n8_w34, c2_n8_w35, c2_n8_w36, c2_n8_w37, c2_n8_w38, c2_n8_w39, c2_n8_w40, c2_n8_w41, c2_n8_w42, c2_n8_w43, c2_n8_w44, c2_n8_w45, c2_n8_w46, c2_n8_w47, c2_n8_w48, c2_n8_w49, c2_n8_w50, c2_n9_w1, c2_n9_w2, c2_n9_w3, c2_n9_w4, c2_n9_w5, c2_n9_w6, c2_n9_w7, c2_n9_w8, c2_n9_w9, c2_n9_w10, c2_n9_w11, c2_n9_w12, c2_n9_w13, c2_n9_w14, c2_n9_w15, c2_n9_w16, c2_n9_w17, c2_n9_w18, c2_n9_w19, c2_n9_w20, c2_n9_w21, c2_n9_w22, c2_n9_w23, c2_n9_w24, c2_n9_w25, c2_n9_w26, c2_n9_w27, c2_n9_w28, c2_n9_w29, c2_n9_w30, c2_n9_w31, c2_n9_w32, c2_n9_w33, c2_n9_w34, c2_n9_w35, c2_n9_w36, c2_n9_w37, c2_n9_w38, c2_n9_w39, c2_n9_w40, c2_n9_w41, c2_n9_w42, c2_n9_w43, c2_n9_w44, c2_n9_w45, c2_n9_w46, c2_n9_w47, c2_n9_w48, c2_n9_w49, c2_n9_w50, c2_n10_w1, c2_n10_w2, c2_n10_w3, c2_n10_w4, c2_n10_w5, c2_n10_w6, c2_n10_w7, c2_n10_w8, c2_n10_w9, c2_n10_w10, c2_n10_w11, c2_n10_w12, c2_n10_w13, c2_n10_w14, c2_n10_w15, c2_n10_w16, c2_n10_w17, c2_n10_w18, c2_n10_w19, c2_n10_w20, c2_n10_w21, c2_n10_w22, c2_n10_w23, c2_n10_w24, c2_n10_w25, c2_n10_w26, c2_n10_w27, c2_n10_w28, c2_n10_w29, c2_n10_w30, c2_n10_w31, c2_n10_w32, c2_n10_w33, c2_n10_w34, c2_n10_w35, c2_n10_w36, c2_n10_w37, c2_n10_w38, c2_n10_w39, c2_n10_w40, c2_n10_w41, c2_n10_w42, c2_n10_w43, c2_n10_w44, c2_n10_w45, c2_n10_w46, c2_n10_w47, c2_n10_w48, c2_n10_w49, c2_n10_w50, c2_n11_w1, c2_n11_w2, c2_n11_w3, c2_n11_w4, c2_n11_w5, c2_n11_w6, c2_n11_w7, c2_n11_w8, c2_n11_w9, c2_n11_w10, c2_n11_w11, c2_n11_w12, c2_n11_w13, c2_n11_w14, c2_n11_w15, c2_n11_w16, c2_n11_w17, c2_n11_w18, c2_n11_w19, c2_n11_w20, c2_n11_w21, c2_n11_w22, c2_n11_w23, c2_n11_w24, c2_n11_w25, c2_n11_w26, c2_n11_w27, c2_n11_w28, c2_n11_w29, c2_n11_w30, c2_n11_w31, c2_n11_w32, c2_n11_w33, c2_n11_w34, c2_n11_w35, c2_n11_w36, c2_n11_w37, c2_n11_w38, c2_n11_w39, c2_n11_w40, c2_n11_w41, c2_n11_w42, c2_n11_w43, c2_n11_w44, c2_n11_w45, c2_n11_w46, c2_n11_w47, c2_n11_w48, c2_n11_w49, c2_n11_w50, c2_n12_w1, c2_n12_w2, c2_n12_w3, c2_n12_w4, c2_n12_w5, c2_n12_w6, c2_n12_w7, c2_n12_w8, c2_n12_w9, c2_n12_w10, c2_n12_w11, c2_n12_w12, c2_n12_w13, c2_n12_w14, c2_n12_w15, c2_n12_w16, c2_n12_w17, c2_n12_w18, c2_n12_w19, c2_n12_w20, c2_n12_w21, c2_n12_w22, c2_n12_w23, c2_n12_w24, c2_n12_w25, c2_n12_w26, c2_n12_w27, c2_n12_w28, c2_n12_w29, c2_n12_w30, c2_n12_w31, c2_n12_w32, c2_n12_w33, c2_n12_w34, c2_n12_w35, c2_n12_w36, c2_n12_w37, c2_n12_w38, c2_n12_w39, c2_n12_w40, c2_n12_w41, c2_n12_w42, c2_n12_w43, c2_n12_w44, c2_n12_w45, c2_n12_w46, c2_n12_w47, c2_n12_w48, c2_n12_w49, c2_n12_w50, c2_n13_w1, c2_n13_w2, c2_n13_w3, c2_n13_w4, c2_n13_w5, c2_n13_w6, c2_n13_w7, c2_n13_w8, c2_n13_w9, c2_n13_w10, c2_n13_w11, c2_n13_w12, c2_n13_w13, c2_n13_w14, c2_n13_w15, c2_n13_w16, c2_n13_w17, c2_n13_w18, c2_n13_w19, c2_n13_w20, c2_n13_w21, c2_n13_w22, c2_n13_w23, c2_n13_w24, c2_n13_w25, c2_n13_w26, c2_n13_w27, c2_n13_w28, c2_n13_w29, c2_n13_w30, c2_n13_w31, c2_n13_w32, c2_n13_w33, c2_n13_w34, c2_n13_w35, c2_n13_w36, c2_n13_w37, c2_n13_w38, c2_n13_w39, c2_n13_w40, c2_n13_w41, c2_n13_w42, c2_n13_w43, c2_n13_w44, c2_n13_w45, c2_n13_w46, c2_n13_w47, c2_n13_w48, c2_n13_w49, c2_n13_w50, c2_n14_w1, c2_n14_w2, c2_n14_w3, c2_n14_w4, c2_n14_w5, c2_n14_w6, c2_n14_w7, c2_n14_w8, c2_n14_w9, c2_n14_w10, c2_n14_w11, c2_n14_w12, c2_n14_w13, c2_n14_w14, c2_n14_w15, c2_n14_w16, c2_n14_w17, c2_n14_w18, c2_n14_w19, c2_n14_w20, c2_n14_w21, c2_n14_w22, c2_n14_w23, c2_n14_w24, c2_n14_w25, c2_n14_w26, c2_n14_w27, c2_n14_w28, c2_n14_w29, c2_n14_w30, c2_n14_w31, c2_n14_w32, c2_n14_w33, c2_n14_w34, c2_n14_w35, c2_n14_w36, c2_n14_w37, c2_n14_w38, c2_n14_w39, c2_n14_w40, c2_n14_w41, c2_n14_w42, c2_n14_w43, c2_n14_w44, c2_n14_w45, c2_n14_w46, c2_n14_w47, c2_n14_w48, c2_n14_w49, c2_n14_w50, c2_n15_w1, c2_n15_w2, c2_n15_w3, c2_n15_w4, c2_n15_w5, c2_n15_w6, c2_n15_w7, c2_n15_w8, c2_n15_w9, c2_n15_w10, c2_n15_w11, c2_n15_w12, c2_n15_w13, c2_n15_w14, c2_n15_w15, c2_n15_w16, c2_n15_w17, c2_n15_w18, c2_n15_w19, c2_n15_w20, c2_n15_w21, c2_n15_w22, c2_n15_w23, c2_n15_w24, c2_n15_w25, c2_n15_w26, c2_n15_w27, c2_n15_w28, c2_n15_w29, c2_n15_w30, c2_n15_w31, c2_n15_w32, c2_n15_w33, c2_n15_w34, c2_n15_w35, c2_n15_w36, c2_n15_w37, c2_n15_w38, c2_n15_w39, c2_n15_w40, c2_n15_w41, c2_n15_w42, c2_n15_w43, c2_n15_w44, c2_n15_w45, c2_n15_w46, c2_n15_w47, c2_n15_w48, c2_n15_w49, c2_n15_w50, c2_n16_w1, c2_n16_w2, c2_n16_w3, c2_n16_w4, c2_n16_w5, c2_n16_w6, c2_n16_w7, c2_n16_w8, c2_n16_w9, c2_n16_w10, c2_n16_w11, c2_n16_w12, c2_n16_w13, c2_n16_w14, c2_n16_w15, c2_n16_w16, c2_n16_w17, c2_n16_w18, c2_n16_w19, c2_n16_w20, c2_n16_w21, c2_n16_w22, c2_n16_w23, c2_n16_w24, c2_n16_w25, c2_n16_w26, c2_n16_w27, c2_n16_w28, c2_n16_w29, c2_n16_w30, c2_n16_w31, c2_n16_w32, c2_n16_w33, c2_n16_w34, c2_n16_w35, c2_n16_w36, c2_n16_w37, c2_n16_w38, c2_n16_w39, c2_n16_w40, c2_n16_w41, c2_n16_w42, c2_n16_w43, c2_n16_w44, c2_n16_w45, c2_n16_w46, c2_n16_w47, c2_n16_w48, c2_n16_w49, c2_n16_w50, c2_n17_w1, c2_n17_w2, c2_n17_w3, c2_n17_w4, c2_n17_w5, c2_n17_w6, c2_n17_w7, c2_n17_w8, c2_n17_w9, c2_n17_w10, c2_n17_w11, c2_n17_w12, c2_n17_w13, c2_n17_w14, c2_n17_w15, c2_n17_w16, c2_n17_w17, c2_n17_w18, c2_n17_w19, c2_n17_w20, c2_n17_w21, c2_n17_w22, c2_n17_w23, c2_n17_w24, c2_n17_w25, c2_n17_w26, c2_n17_w27, c2_n17_w28, c2_n17_w29, c2_n17_w30, c2_n17_w31, c2_n17_w32, c2_n17_w33, c2_n17_w34, c2_n17_w35, c2_n17_w36, c2_n17_w37, c2_n17_w38, c2_n17_w39, c2_n17_w40, c2_n17_w41, c2_n17_w42, c2_n17_w43, c2_n17_w44, c2_n17_w45, c2_n17_w46, c2_n17_w47, c2_n17_w48, c2_n17_w49, c2_n17_w50, c2_n18_w1, c2_n18_w2, c2_n18_w3, c2_n18_w4, c2_n18_w5, c2_n18_w6, c2_n18_w7, c2_n18_w8, c2_n18_w9, c2_n18_w10, c2_n18_w11, c2_n18_w12, c2_n18_w13, c2_n18_w14, c2_n18_w15, c2_n18_w16, c2_n18_w17, c2_n18_w18, c2_n18_w19, c2_n18_w20, c2_n18_w21, c2_n18_w22, c2_n18_w23, c2_n18_w24, c2_n18_w25, c2_n18_w26, c2_n18_w27, c2_n18_w28, c2_n18_w29, c2_n18_w30, c2_n18_w31, c2_n18_w32, c2_n18_w33, c2_n18_w34, c2_n18_w35, c2_n18_w36, c2_n18_w37, c2_n18_w38, c2_n18_w39, c2_n18_w40, c2_n18_w41, c2_n18_w42, c2_n18_w43, c2_n18_w44, c2_n18_w45, c2_n18_w46, c2_n18_w47, c2_n18_w48, c2_n18_w49, c2_n18_w50, c2_n19_w1, c2_n19_w2, c2_n19_w3, c2_n19_w4, c2_n19_w5, c2_n19_w6, c2_n19_w7, c2_n19_w8, c2_n19_w9, c2_n19_w10, c2_n19_w11, c2_n19_w12, c2_n19_w13, c2_n19_w14, c2_n19_w15, c2_n19_w16, c2_n19_w17, c2_n19_w18, c2_n19_w19, c2_n19_w20, c2_n19_w21, c2_n19_w22, c2_n19_w23, c2_n19_w24, c2_n19_w25, c2_n19_w26, c2_n19_w27, c2_n19_w28, c2_n19_w29, c2_n19_w30, c2_n19_w31, c2_n19_w32, c2_n19_w33, c2_n19_w34, c2_n19_w35, c2_n19_w36, c2_n19_w37, c2_n19_w38, c2_n19_w39, c2_n19_w40, c2_n19_w41, c2_n19_w42, c2_n19_w43, c2_n19_w44, c2_n19_w45, c2_n19_w46, c2_n19_w47, c2_n19_w48, c2_n19_w49, c2_n19_w50, c2_n20_w1, c2_n20_w2, c2_n20_w3, c2_n20_w4, c2_n20_w5, c2_n20_w6, c2_n20_w7, c2_n20_w8, c2_n20_w9, c2_n20_w10, c2_n20_w11, c2_n20_w12, c2_n20_w13, c2_n20_w14, c2_n20_w15, c2_n20_w16, c2_n20_w17, c2_n20_w18, c2_n20_w19, c2_n20_w20, c2_n20_w21, c2_n20_w22, c2_n20_w23, c2_n20_w24, c2_n20_w25, c2_n20_w26, c2_n20_w27, c2_n20_w28, c2_n20_w29, c2_n20_w30, c2_n20_w31, c2_n20_w32, c2_n20_w33, c2_n20_w34, c2_n20_w35, c2_n20_w36, c2_n20_w37, c2_n20_w38, c2_n20_w39, c2_n20_w40, c2_n20_w41, c2_n20_w42, c2_n20_w43, c2_n20_w44, c2_n20_w45, c2_n20_w46, c2_n20_w47, c2_n20_w48, c2_n20_w49, c2_n20_w50, c2_n21_w1, c2_n21_w2, c2_n21_w3, c2_n21_w4, c2_n21_w5, c2_n21_w6, c2_n21_w7, c2_n21_w8, c2_n21_w9, c2_n21_w10, c2_n21_w11, c2_n21_w12, c2_n21_w13, c2_n21_w14, c2_n21_w15, c2_n21_w16, c2_n21_w17, c2_n21_w18, c2_n21_w19, c2_n21_w20, c2_n21_w21, c2_n21_w22, c2_n21_w23, c2_n21_w24, c2_n21_w25, c2_n21_w26, c2_n21_w27, c2_n21_w28, c2_n21_w29, c2_n21_w30, c2_n21_w31, c2_n21_w32, c2_n21_w33, c2_n21_w34, c2_n21_w35, c2_n21_w36, c2_n21_w37, c2_n21_w38, c2_n21_w39, c2_n21_w40, c2_n21_w41, c2_n21_w42, c2_n21_w43, c2_n21_w44, c2_n21_w45, c2_n21_w46, c2_n21_w47, c2_n21_w48, c2_n21_w49, c2_n21_w50, c2_n22_w1, c2_n22_w2, c2_n22_w3, c2_n22_w4, c2_n22_w5, c2_n22_w6, c2_n22_w7, c2_n22_w8, c2_n22_w9, c2_n22_w10, c2_n22_w11, c2_n22_w12, c2_n22_w13, c2_n22_w14, c2_n22_w15, c2_n22_w16, c2_n22_w17, c2_n22_w18, c2_n22_w19, c2_n22_w20, c2_n22_w21, c2_n22_w22, c2_n22_w23, c2_n22_w24, c2_n22_w25, c2_n22_w26, c2_n22_w27, c2_n22_w28, c2_n22_w29, c2_n22_w30, c2_n22_w31, c2_n22_w32, c2_n22_w33, c2_n22_w34, c2_n22_w35, c2_n22_w36, c2_n22_w37, c2_n22_w38, c2_n22_w39, c2_n22_w40, c2_n22_w41, c2_n22_w42, c2_n22_w43, c2_n22_w44, c2_n22_w45, c2_n22_w46, c2_n22_w47, c2_n22_w48, c2_n22_w49, c2_n22_w50, c2_n23_w1, c2_n23_w2, c2_n23_w3, c2_n23_w4, c2_n23_w5, c2_n23_w6, c2_n23_w7, c2_n23_w8, c2_n23_w9, c2_n23_w10, c2_n23_w11, c2_n23_w12, c2_n23_w13, c2_n23_w14, c2_n23_w15, c2_n23_w16, c2_n23_w17, c2_n23_w18, c2_n23_w19, c2_n23_w20, c2_n23_w21, c2_n23_w22, c2_n23_w23, c2_n23_w24, c2_n23_w25, c2_n23_w26, c2_n23_w27, c2_n23_w28, c2_n23_w29, c2_n23_w30, c2_n23_w31, c2_n23_w32, c2_n23_w33, c2_n23_w34, c2_n23_w35, c2_n23_w36, c2_n23_w37, c2_n23_w38, c2_n23_w39, c2_n23_w40, c2_n23_w41, c2_n23_w42, c2_n23_w43, c2_n23_w44, c2_n23_w45, c2_n23_w46, c2_n23_w47, c2_n23_w48, c2_n23_w49, c2_n23_w50, c2_n24_w1, c2_n24_w2, c2_n24_w3, c2_n24_w4, c2_n24_w5, c2_n24_w6, c2_n24_w7, c2_n24_w8, c2_n24_w9, c2_n24_w10, c2_n24_w11, c2_n24_w12, c2_n24_w13, c2_n24_w14, c2_n24_w15, c2_n24_w16, c2_n24_w17, c2_n24_w18, c2_n24_w19, c2_n24_w20, c2_n24_w21, c2_n24_w22, c2_n24_w23, c2_n24_w24, c2_n24_w25, c2_n24_w26, c2_n24_w27, c2_n24_w28, c2_n24_w29, c2_n24_w30, c2_n24_w31, c2_n24_w32, c2_n24_w33, c2_n24_w34, c2_n24_w35, c2_n24_w36, c2_n24_w37, c2_n24_w38, c2_n24_w39, c2_n24_w40, c2_n24_w41, c2_n24_w42, c2_n24_w43, c2_n24_w44, c2_n24_w45, c2_n24_w46, c2_n24_w47, c2_n24_w48, c2_n24_w49, c2_n24_w50, c2_n25_w1, c2_n25_w2, c2_n25_w3, c2_n25_w4, c2_n25_w5, c2_n25_w6, c2_n25_w7, c2_n25_w8, c2_n25_w9, c2_n25_w10, c2_n25_w11, c2_n25_w12, c2_n25_w13, c2_n25_w14, c2_n25_w15, c2_n25_w16, c2_n25_w17, c2_n25_w18, c2_n25_w19, c2_n25_w20, c2_n25_w21, c2_n25_w22, c2_n25_w23, c2_n25_w24, c2_n25_w25, c2_n25_w26, c2_n25_w27, c2_n25_w28, c2_n25_w29, c2_n25_w30, c2_n25_w31, c2_n25_w32, c2_n25_w33, c2_n25_w34, c2_n25_w35, c2_n25_w36, c2_n25_w37, c2_n25_w38, c2_n25_w39, c2_n25_w40, c2_n25_w41, c2_n25_w42, c2_n25_w43, c2_n25_w44, c2_n25_w45, c2_n25_w46, c2_n25_w47, c2_n25_w48, c2_n25_w49, c2_n25_w50, c2_n26_w1, c2_n26_w2, c2_n26_w3, c2_n26_w4, c2_n26_w5, c2_n26_w6, c2_n26_w7, c2_n26_w8, c2_n26_w9, c2_n26_w10, c2_n26_w11, c2_n26_w12, c2_n26_w13, c2_n26_w14, c2_n26_w15, c2_n26_w16, c2_n26_w17, c2_n26_w18, c2_n26_w19, c2_n26_w20, c2_n26_w21, c2_n26_w22, c2_n26_w23, c2_n26_w24, c2_n26_w25, c2_n26_w26, c2_n26_w27, c2_n26_w28, c2_n26_w29, c2_n26_w30, c2_n26_w31, c2_n26_w32, c2_n26_w33, c2_n26_w34, c2_n26_w35, c2_n26_w36, c2_n26_w37, c2_n26_w38, c2_n26_w39, c2_n26_w40, c2_n26_w41, c2_n26_w42, c2_n26_w43, c2_n26_w44, c2_n26_w45, c2_n26_w46, c2_n26_w47, c2_n26_w48, c2_n26_w49, c2_n26_w50, c2_n27_w1, c2_n27_w2, c2_n27_w3, c2_n27_w4, c2_n27_w5, c2_n27_w6, c2_n27_w7, c2_n27_w8, c2_n27_w9, c2_n27_w10, c2_n27_w11, c2_n27_w12, c2_n27_w13, c2_n27_w14, c2_n27_w15, c2_n27_w16, c2_n27_w17, c2_n27_w18, c2_n27_w19, c2_n27_w20, c2_n27_w21, c2_n27_w22, c2_n27_w23, c2_n27_w24, c2_n27_w25, c2_n27_w26, c2_n27_w27, c2_n27_w28, c2_n27_w29, c2_n27_w30, c2_n27_w31, c2_n27_w32, c2_n27_w33, c2_n27_w34, c2_n27_w35, c2_n27_w36, c2_n27_w37, c2_n27_w38, c2_n27_w39, c2_n27_w40, c2_n27_w41, c2_n27_w42, c2_n27_w43, c2_n27_w44, c2_n27_w45, c2_n27_w46, c2_n27_w47, c2_n27_w48, c2_n27_w49, c2_n27_w50, c2_n28_w1, c2_n28_w2, c2_n28_w3, c2_n28_w4, c2_n28_w5, c2_n28_w6, c2_n28_w7, c2_n28_w8, c2_n28_w9, c2_n28_w10, c2_n28_w11, c2_n28_w12, c2_n28_w13, c2_n28_w14, c2_n28_w15, c2_n28_w16, c2_n28_w17, c2_n28_w18, c2_n28_w19, c2_n28_w20, c2_n28_w21, c2_n28_w22, c2_n28_w23, c2_n28_w24, c2_n28_w25, c2_n28_w26, c2_n28_w27, c2_n28_w28, c2_n28_w29, c2_n28_w30, c2_n28_w31, c2_n28_w32, c2_n28_w33, c2_n28_w34, c2_n28_w35, c2_n28_w36, c2_n28_w37, c2_n28_w38, c2_n28_w39, c2_n28_w40, c2_n28_w41, c2_n28_w42, c2_n28_w43, c2_n28_w44, c2_n28_w45, c2_n28_w46, c2_n28_w47, c2_n28_w48, c2_n28_w49, c2_n28_w50, c2_n29_w1, c2_n29_w2, c2_n29_w3, c2_n29_w4, c2_n29_w5, c2_n29_w6, c2_n29_w7, c2_n29_w8, c2_n29_w9, c2_n29_w10, c2_n29_w11, c2_n29_w12, c2_n29_w13, c2_n29_w14, c2_n29_w15, c2_n29_w16, c2_n29_w17, c2_n29_w18, c2_n29_w19, c2_n29_w20, c2_n29_w21, c2_n29_w22, c2_n29_w23, c2_n29_w24, c2_n29_w25, c2_n29_w26, c2_n29_w27, c2_n29_w28, c2_n29_w29, c2_n29_w30, c2_n29_w31, c2_n29_w32, c2_n29_w33, c2_n29_w34, c2_n29_w35, c2_n29_w36, c2_n29_w37, c2_n29_w38, c2_n29_w39, c2_n29_w40, c2_n29_w41, c2_n29_w42, c2_n29_w43, c2_n29_w44, c2_n29_w45, c2_n29_w46, c2_n29_w47, c2_n29_w48, c2_n29_w49, c2_n29_w50: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c2_n0_y, c2_n1_y, c2_n2_y, c2_n3_y, c2_n4_y, c2_n5_y, c2_n6_y, c2_n7_y, c2_n8_y, c2_n9_y, c2_n10_y, c2_n11_y, c2_n12_y, c2_n13_y, c2_n14_y, c2_n15_y, c2_n16_y, c2_n17_y, c2_n18_y, c2_n19_y, c2_n20_y, c2_n21_y, c2_n22_y, c2_n23_y, c2_n24_y, c2_n25_y, c2_n26_y, c2_n27_y, c2_n28_y, c2_n29_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada2_ReLU_30neuron_8bits_50n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n0_w1, 
            w2=> c2_n0_w2, 
            w3=> c2_n0_w3, 
            w4=> c2_n0_w4, 
            w5=> c2_n0_w5, 
            w6=> c2_n0_w6, 
            w7=> c2_n0_w7, 
            w8=> c2_n0_w8, 
            w9=> c2_n0_w9, 
            w10=> c2_n0_w10, 
            w11=> c2_n0_w11, 
            w12=> c2_n0_w12, 
            w13=> c2_n0_w13, 
            w14=> c2_n0_w14, 
            w15=> c2_n0_w15, 
            w16=> c2_n0_w16, 
            w17=> c2_n0_w17, 
            w18=> c2_n0_w18, 
            w19=> c2_n0_w19, 
            w20=> c2_n0_w20, 
            w21=> c2_n0_w21, 
            w22=> c2_n0_w22, 
            w23=> c2_n0_w23, 
            w24=> c2_n0_w24, 
            w25=> c2_n0_w25, 
            w26=> c2_n0_w26, 
            w27=> c2_n0_w27, 
            w28=> c2_n0_w28, 
            w29=> c2_n0_w29, 
            w30=> c2_n0_w30, 
            w31=> c2_n0_w31, 
            w32=> c2_n0_w32, 
            w33=> c2_n0_w33, 
            w34=> c2_n0_w34, 
            w35=> c2_n0_w35, 
            w36=> c2_n0_w36, 
            w37=> c2_n0_w37, 
            w38=> c2_n0_w38, 
            w39=> c2_n0_w39, 
            w40=> c2_n0_w40, 
            w41=> c2_n0_w41, 
            w42=> c2_n0_w42, 
            w43=> c2_n0_w43, 
            w44=> c2_n0_w44, 
            w45=> c2_n0_w45, 
            w46=> c2_n0_w46, 
            w47=> c2_n0_w47, 
            w48=> c2_n0_w48, 
            w49=> c2_n0_w49, 
            w50=> c2_n0_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n1_w1, 
            w2=> c2_n1_w2, 
            w3=> c2_n1_w3, 
            w4=> c2_n1_w4, 
            w5=> c2_n1_w5, 
            w6=> c2_n1_w6, 
            w7=> c2_n1_w7, 
            w8=> c2_n1_w8, 
            w9=> c2_n1_w9, 
            w10=> c2_n1_w10, 
            w11=> c2_n1_w11, 
            w12=> c2_n1_w12, 
            w13=> c2_n1_w13, 
            w14=> c2_n1_w14, 
            w15=> c2_n1_w15, 
            w16=> c2_n1_w16, 
            w17=> c2_n1_w17, 
            w18=> c2_n1_w18, 
            w19=> c2_n1_w19, 
            w20=> c2_n1_w20, 
            w21=> c2_n1_w21, 
            w22=> c2_n1_w22, 
            w23=> c2_n1_w23, 
            w24=> c2_n1_w24, 
            w25=> c2_n1_w25, 
            w26=> c2_n1_w26, 
            w27=> c2_n1_w27, 
            w28=> c2_n1_w28, 
            w29=> c2_n1_w29, 
            w30=> c2_n1_w30, 
            w31=> c2_n1_w31, 
            w32=> c2_n1_w32, 
            w33=> c2_n1_w33, 
            w34=> c2_n1_w34, 
            w35=> c2_n1_w35, 
            w36=> c2_n1_w36, 
            w37=> c2_n1_w37, 
            w38=> c2_n1_w38, 
            w39=> c2_n1_w39, 
            w40=> c2_n1_w40, 
            w41=> c2_n1_w41, 
            w42=> c2_n1_w42, 
            w43=> c2_n1_w43, 
            w44=> c2_n1_w44, 
            w45=> c2_n1_w45, 
            w46=> c2_n1_w46, 
            w47=> c2_n1_w47, 
            w48=> c2_n1_w48, 
            w49=> c2_n1_w49, 
            w50=> c2_n1_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n2_w1, 
            w2=> c2_n2_w2, 
            w3=> c2_n2_w3, 
            w4=> c2_n2_w4, 
            w5=> c2_n2_w5, 
            w6=> c2_n2_w6, 
            w7=> c2_n2_w7, 
            w8=> c2_n2_w8, 
            w9=> c2_n2_w9, 
            w10=> c2_n2_w10, 
            w11=> c2_n2_w11, 
            w12=> c2_n2_w12, 
            w13=> c2_n2_w13, 
            w14=> c2_n2_w14, 
            w15=> c2_n2_w15, 
            w16=> c2_n2_w16, 
            w17=> c2_n2_w17, 
            w18=> c2_n2_w18, 
            w19=> c2_n2_w19, 
            w20=> c2_n2_w20, 
            w21=> c2_n2_w21, 
            w22=> c2_n2_w22, 
            w23=> c2_n2_w23, 
            w24=> c2_n2_w24, 
            w25=> c2_n2_w25, 
            w26=> c2_n2_w26, 
            w27=> c2_n2_w27, 
            w28=> c2_n2_w28, 
            w29=> c2_n2_w29, 
            w30=> c2_n2_w30, 
            w31=> c2_n2_w31, 
            w32=> c2_n2_w32, 
            w33=> c2_n2_w33, 
            w34=> c2_n2_w34, 
            w35=> c2_n2_w35, 
            w36=> c2_n2_w36, 
            w37=> c2_n2_w37, 
            w38=> c2_n2_w38, 
            w39=> c2_n2_w39, 
            w40=> c2_n2_w40, 
            w41=> c2_n2_w41, 
            w42=> c2_n2_w42, 
            w43=> c2_n2_w43, 
            w44=> c2_n2_w44, 
            w45=> c2_n2_w45, 
            w46=> c2_n2_w46, 
            w47=> c2_n2_w47, 
            w48=> c2_n2_w48, 
            w49=> c2_n2_w49, 
            w50=> c2_n2_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n3_w1, 
            w2=> c2_n3_w2, 
            w3=> c2_n3_w3, 
            w4=> c2_n3_w4, 
            w5=> c2_n3_w5, 
            w6=> c2_n3_w6, 
            w7=> c2_n3_w7, 
            w8=> c2_n3_w8, 
            w9=> c2_n3_w9, 
            w10=> c2_n3_w10, 
            w11=> c2_n3_w11, 
            w12=> c2_n3_w12, 
            w13=> c2_n3_w13, 
            w14=> c2_n3_w14, 
            w15=> c2_n3_w15, 
            w16=> c2_n3_w16, 
            w17=> c2_n3_w17, 
            w18=> c2_n3_w18, 
            w19=> c2_n3_w19, 
            w20=> c2_n3_w20, 
            w21=> c2_n3_w21, 
            w22=> c2_n3_w22, 
            w23=> c2_n3_w23, 
            w24=> c2_n3_w24, 
            w25=> c2_n3_w25, 
            w26=> c2_n3_w26, 
            w27=> c2_n3_w27, 
            w28=> c2_n3_w28, 
            w29=> c2_n3_w29, 
            w30=> c2_n3_w30, 
            w31=> c2_n3_w31, 
            w32=> c2_n3_w32, 
            w33=> c2_n3_w33, 
            w34=> c2_n3_w34, 
            w35=> c2_n3_w35, 
            w36=> c2_n3_w36, 
            w37=> c2_n3_w37, 
            w38=> c2_n3_w38, 
            w39=> c2_n3_w39, 
            w40=> c2_n3_w40, 
            w41=> c2_n3_w41, 
            w42=> c2_n3_w42, 
            w43=> c2_n3_w43, 
            w44=> c2_n3_w44, 
            w45=> c2_n3_w45, 
            w46=> c2_n3_w46, 
            w47=> c2_n3_w47, 
            w48=> c2_n3_w48, 
            w49=> c2_n3_w49, 
            w50=> c2_n3_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n4_w1, 
            w2=> c2_n4_w2, 
            w3=> c2_n4_w3, 
            w4=> c2_n4_w4, 
            w5=> c2_n4_w5, 
            w6=> c2_n4_w6, 
            w7=> c2_n4_w7, 
            w8=> c2_n4_w8, 
            w9=> c2_n4_w9, 
            w10=> c2_n4_w10, 
            w11=> c2_n4_w11, 
            w12=> c2_n4_w12, 
            w13=> c2_n4_w13, 
            w14=> c2_n4_w14, 
            w15=> c2_n4_w15, 
            w16=> c2_n4_w16, 
            w17=> c2_n4_w17, 
            w18=> c2_n4_w18, 
            w19=> c2_n4_w19, 
            w20=> c2_n4_w20, 
            w21=> c2_n4_w21, 
            w22=> c2_n4_w22, 
            w23=> c2_n4_w23, 
            w24=> c2_n4_w24, 
            w25=> c2_n4_w25, 
            w26=> c2_n4_w26, 
            w27=> c2_n4_w27, 
            w28=> c2_n4_w28, 
            w29=> c2_n4_w29, 
            w30=> c2_n4_w30, 
            w31=> c2_n4_w31, 
            w32=> c2_n4_w32, 
            w33=> c2_n4_w33, 
            w34=> c2_n4_w34, 
            w35=> c2_n4_w35, 
            w36=> c2_n4_w36, 
            w37=> c2_n4_w37, 
            w38=> c2_n4_w38, 
            w39=> c2_n4_w39, 
            w40=> c2_n4_w40, 
            w41=> c2_n4_w41, 
            w42=> c2_n4_w42, 
            w43=> c2_n4_w43, 
            w44=> c2_n4_w44, 
            w45=> c2_n4_w45, 
            w46=> c2_n4_w46, 
            w47=> c2_n4_w47, 
            w48=> c2_n4_w48, 
            w49=> c2_n4_w49, 
            w50=> c2_n4_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n5_w1, 
            w2=> c2_n5_w2, 
            w3=> c2_n5_w3, 
            w4=> c2_n5_w4, 
            w5=> c2_n5_w5, 
            w6=> c2_n5_w6, 
            w7=> c2_n5_w7, 
            w8=> c2_n5_w8, 
            w9=> c2_n5_w9, 
            w10=> c2_n5_w10, 
            w11=> c2_n5_w11, 
            w12=> c2_n5_w12, 
            w13=> c2_n5_w13, 
            w14=> c2_n5_w14, 
            w15=> c2_n5_w15, 
            w16=> c2_n5_w16, 
            w17=> c2_n5_w17, 
            w18=> c2_n5_w18, 
            w19=> c2_n5_w19, 
            w20=> c2_n5_w20, 
            w21=> c2_n5_w21, 
            w22=> c2_n5_w22, 
            w23=> c2_n5_w23, 
            w24=> c2_n5_w24, 
            w25=> c2_n5_w25, 
            w26=> c2_n5_w26, 
            w27=> c2_n5_w27, 
            w28=> c2_n5_w28, 
            w29=> c2_n5_w29, 
            w30=> c2_n5_w30, 
            w31=> c2_n5_w31, 
            w32=> c2_n5_w32, 
            w33=> c2_n5_w33, 
            w34=> c2_n5_w34, 
            w35=> c2_n5_w35, 
            w36=> c2_n5_w36, 
            w37=> c2_n5_w37, 
            w38=> c2_n5_w38, 
            w39=> c2_n5_w39, 
            w40=> c2_n5_w40, 
            w41=> c2_n5_w41, 
            w42=> c2_n5_w42, 
            w43=> c2_n5_w43, 
            w44=> c2_n5_w44, 
            w45=> c2_n5_w45, 
            w46=> c2_n5_w46, 
            w47=> c2_n5_w47, 
            w48=> c2_n5_w48, 
            w49=> c2_n5_w49, 
            w50=> c2_n5_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n6_w1, 
            w2=> c2_n6_w2, 
            w3=> c2_n6_w3, 
            w4=> c2_n6_w4, 
            w5=> c2_n6_w5, 
            w6=> c2_n6_w6, 
            w7=> c2_n6_w7, 
            w8=> c2_n6_w8, 
            w9=> c2_n6_w9, 
            w10=> c2_n6_w10, 
            w11=> c2_n6_w11, 
            w12=> c2_n6_w12, 
            w13=> c2_n6_w13, 
            w14=> c2_n6_w14, 
            w15=> c2_n6_w15, 
            w16=> c2_n6_w16, 
            w17=> c2_n6_w17, 
            w18=> c2_n6_w18, 
            w19=> c2_n6_w19, 
            w20=> c2_n6_w20, 
            w21=> c2_n6_w21, 
            w22=> c2_n6_w22, 
            w23=> c2_n6_w23, 
            w24=> c2_n6_w24, 
            w25=> c2_n6_w25, 
            w26=> c2_n6_w26, 
            w27=> c2_n6_w27, 
            w28=> c2_n6_w28, 
            w29=> c2_n6_w29, 
            w30=> c2_n6_w30, 
            w31=> c2_n6_w31, 
            w32=> c2_n6_w32, 
            w33=> c2_n6_w33, 
            w34=> c2_n6_w34, 
            w35=> c2_n6_w35, 
            w36=> c2_n6_w36, 
            w37=> c2_n6_w37, 
            w38=> c2_n6_w38, 
            w39=> c2_n6_w39, 
            w40=> c2_n6_w40, 
            w41=> c2_n6_w41, 
            w42=> c2_n6_w42, 
            w43=> c2_n6_w43, 
            w44=> c2_n6_w44, 
            w45=> c2_n6_w45, 
            w46=> c2_n6_w46, 
            w47=> c2_n6_w47, 
            w48=> c2_n6_w48, 
            w49=> c2_n6_w49, 
            w50=> c2_n6_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n7_w1, 
            w2=> c2_n7_w2, 
            w3=> c2_n7_w3, 
            w4=> c2_n7_w4, 
            w5=> c2_n7_w5, 
            w6=> c2_n7_w6, 
            w7=> c2_n7_w7, 
            w8=> c2_n7_w8, 
            w9=> c2_n7_w9, 
            w10=> c2_n7_w10, 
            w11=> c2_n7_w11, 
            w12=> c2_n7_w12, 
            w13=> c2_n7_w13, 
            w14=> c2_n7_w14, 
            w15=> c2_n7_w15, 
            w16=> c2_n7_w16, 
            w17=> c2_n7_w17, 
            w18=> c2_n7_w18, 
            w19=> c2_n7_w19, 
            w20=> c2_n7_w20, 
            w21=> c2_n7_w21, 
            w22=> c2_n7_w22, 
            w23=> c2_n7_w23, 
            w24=> c2_n7_w24, 
            w25=> c2_n7_w25, 
            w26=> c2_n7_w26, 
            w27=> c2_n7_w27, 
            w28=> c2_n7_w28, 
            w29=> c2_n7_w29, 
            w30=> c2_n7_w30, 
            w31=> c2_n7_w31, 
            w32=> c2_n7_w32, 
            w33=> c2_n7_w33, 
            w34=> c2_n7_w34, 
            w35=> c2_n7_w35, 
            w36=> c2_n7_w36, 
            w37=> c2_n7_w37, 
            w38=> c2_n7_w38, 
            w39=> c2_n7_w39, 
            w40=> c2_n7_w40, 
            w41=> c2_n7_w41, 
            w42=> c2_n7_w42, 
            w43=> c2_n7_w43, 
            w44=> c2_n7_w44, 
            w45=> c2_n7_w45, 
            w46=> c2_n7_w46, 
            w47=> c2_n7_w47, 
            w48=> c2_n7_w48, 
            w49=> c2_n7_w49, 
            w50=> c2_n7_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n8_w1, 
            w2=> c2_n8_w2, 
            w3=> c2_n8_w3, 
            w4=> c2_n8_w4, 
            w5=> c2_n8_w5, 
            w6=> c2_n8_w6, 
            w7=> c2_n8_w7, 
            w8=> c2_n8_w8, 
            w9=> c2_n8_w9, 
            w10=> c2_n8_w10, 
            w11=> c2_n8_w11, 
            w12=> c2_n8_w12, 
            w13=> c2_n8_w13, 
            w14=> c2_n8_w14, 
            w15=> c2_n8_w15, 
            w16=> c2_n8_w16, 
            w17=> c2_n8_w17, 
            w18=> c2_n8_w18, 
            w19=> c2_n8_w19, 
            w20=> c2_n8_w20, 
            w21=> c2_n8_w21, 
            w22=> c2_n8_w22, 
            w23=> c2_n8_w23, 
            w24=> c2_n8_w24, 
            w25=> c2_n8_w25, 
            w26=> c2_n8_w26, 
            w27=> c2_n8_w27, 
            w28=> c2_n8_w28, 
            w29=> c2_n8_w29, 
            w30=> c2_n8_w30, 
            w31=> c2_n8_w31, 
            w32=> c2_n8_w32, 
            w33=> c2_n8_w33, 
            w34=> c2_n8_w34, 
            w35=> c2_n8_w35, 
            w36=> c2_n8_w36, 
            w37=> c2_n8_w37, 
            w38=> c2_n8_w38, 
            w39=> c2_n8_w39, 
            w40=> c2_n8_w40, 
            w41=> c2_n8_w41, 
            w42=> c2_n8_w42, 
            w43=> c2_n8_w43, 
            w44=> c2_n8_w44, 
            w45=> c2_n8_w45, 
            w46=> c2_n8_w46, 
            w47=> c2_n8_w47, 
            w48=> c2_n8_w48, 
            w49=> c2_n8_w49, 
            w50=> c2_n8_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n9_w1, 
            w2=> c2_n9_w2, 
            w3=> c2_n9_w3, 
            w4=> c2_n9_w4, 
            w5=> c2_n9_w5, 
            w6=> c2_n9_w6, 
            w7=> c2_n9_w7, 
            w8=> c2_n9_w8, 
            w9=> c2_n9_w9, 
            w10=> c2_n9_w10, 
            w11=> c2_n9_w11, 
            w12=> c2_n9_w12, 
            w13=> c2_n9_w13, 
            w14=> c2_n9_w14, 
            w15=> c2_n9_w15, 
            w16=> c2_n9_w16, 
            w17=> c2_n9_w17, 
            w18=> c2_n9_w18, 
            w19=> c2_n9_w19, 
            w20=> c2_n9_w20, 
            w21=> c2_n9_w21, 
            w22=> c2_n9_w22, 
            w23=> c2_n9_w23, 
            w24=> c2_n9_w24, 
            w25=> c2_n9_w25, 
            w26=> c2_n9_w26, 
            w27=> c2_n9_w27, 
            w28=> c2_n9_w28, 
            w29=> c2_n9_w29, 
            w30=> c2_n9_w30, 
            w31=> c2_n9_w31, 
            w32=> c2_n9_w32, 
            w33=> c2_n9_w33, 
            w34=> c2_n9_w34, 
            w35=> c2_n9_w35, 
            w36=> c2_n9_w36, 
            w37=> c2_n9_w37, 
            w38=> c2_n9_w38, 
            w39=> c2_n9_w39, 
            w40=> c2_n9_w40, 
            w41=> c2_n9_w41, 
            w42=> c2_n9_w42, 
            w43=> c2_n9_w43, 
            w44=> c2_n9_w44, 
            w45=> c2_n9_w45, 
            w46=> c2_n9_w46, 
            w47=> c2_n9_w47, 
            w48=> c2_n9_w48, 
            w49=> c2_n9_w49, 
            w50=> c2_n9_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n9_y
   );           
            
neuron_inst_10: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n10_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n10_w1, 
            w2=> c2_n10_w2, 
            w3=> c2_n10_w3, 
            w4=> c2_n10_w4, 
            w5=> c2_n10_w5, 
            w6=> c2_n10_w6, 
            w7=> c2_n10_w7, 
            w8=> c2_n10_w8, 
            w9=> c2_n10_w9, 
            w10=> c2_n10_w10, 
            w11=> c2_n10_w11, 
            w12=> c2_n10_w12, 
            w13=> c2_n10_w13, 
            w14=> c2_n10_w14, 
            w15=> c2_n10_w15, 
            w16=> c2_n10_w16, 
            w17=> c2_n10_w17, 
            w18=> c2_n10_w18, 
            w19=> c2_n10_w19, 
            w20=> c2_n10_w20, 
            w21=> c2_n10_w21, 
            w22=> c2_n10_w22, 
            w23=> c2_n10_w23, 
            w24=> c2_n10_w24, 
            w25=> c2_n10_w25, 
            w26=> c2_n10_w26, 
            w27=> c2_n10_w27, 
            w28=> c2_n10_w28, 
            w29=> c2_n10_w29, 
            w30=> c2_n10_w30, 
            w31=> c2_n10_w31, 
            w32=> c2_n10_w32, 
            w33=> c2_n10_w33, 
            w34=> c2_n10_w34, 
            w35=> c2_n10_w35, 
            w36=> c2_n10_w36, 
            w37=> c2_n10_w37, 
            w38=> c2_n10_w38, 
            w39=> c2_n10_w39, 
            w40=> c2_n10_w40, 
            w41=> c2_n10_w41, 
            w42=> c2_n10_w42, 
            w43=> c2_n10_w43, 
            w44=> c2_n10_w44, 
            w45=> c2_n10_w45, 
            w46=> c2_n10_w46, 
            w47=> c2_n10_w47, 
            w48=> c2_n10_w48, 
            w49=> c2_n10_w49, 
            w50=> c2_n10_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n10_y
   );           
            
neuron_inst_11: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n11_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n11_w1, 
            w2=> c2_n11_w2, 
            w3=> c2_n11_w3, 
            w4=> c2_n11_w4, 
            w5=> c2_n11_w5, 
            w6=> c2_n11_w6, 
            w7=> c2_n11_w7, 
            w8=> c2_n11_w8, 
            w9=> c2_n11_w9, 
            w10=> c2_n11_w10, 
            w11=> c2_n11_w11, 
            w12=> c2_n11_w12, 
            w13=> c2_n11_w13, 
            w14=> c2_n11_w14, 
            w15=> c2_n11_w15, 
            w16=> c2_n11_w16, 
            w17=> c2_n11_w17, 
            w18=> c2_n11_w18, 
            w19=> c2_n11_w19, 
            w20=> c2_n11_w20, 
            w21=> c2_n11_w21, 
            w22=> c2_n11_w22, 
            w23=> c2_n11_w23, 
            w24=> c2_n11_w24, 
            w25=> c2_n11_w25, 
            w26=> c2_n11_w26, 
            w27=> c2_n11_w27, 
            w28=> c2_n11_w28, 
            w29=> c2_n11_w29, 
            w30=> c2_n11_w30, 
            w31=> c2_n11_w31, 
            w32=> c2_n11_w32, 
            w33=> c2_n11_w33, 
            w34=> c2_n11_w34, 
            w35=> c2_n11_w35, 
            w36=> c2_n11_w36, 
            w37=> c2_n11_w37, 
            w38=> c2_n11_w38, 
            w39=> c2_n11_w39, 
            w40=> c2_n11_w40, 
            w41=> c2_n11_w41, 
            w42=> c2_n11_w42, 
            w43=> c2_n11_w43, 
            w44=> c2_n11_w44, 
            w45=> c2_n11_w45, 
            w46=> c2_n11_w46, 
            w47=> c2_n11_w47, 
            w48=> c2_n11_w48, 
            w49=> c2_n11_w49, 
            w50=> c2_n11_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n11_y
   );           
            
neuron_inst_12: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n12_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n12_w1, 
            w2=> c2_n12_w2, 
            w3=> c2_n12_w3, 
            w4=> c2_n12_w4, 
            w5=> c2_n12_w5, 
            w6=> c2_n12_w6, 
            w7=> c2_n12_w7, 
            w8=> c2_n12_w8, 
            w9=> c2_n12_w9, 
            w10=> c2_n12_w10, 
            w11=> c2_n12_w11, 
            w12=> c2_n12_w12, 
            w13=> c2_n12_w13, 
            w14=> c2_n12_w14, 
            w15=> c2_n12_w15, 
            w16=> c2_n12_w16, 
            w17=> c2_n12_w17, 
            w18=> c2_n12_w18, 
            w19=> c2_n12_w19, 
            w20=> c2_n12_w20, 
            w21=> c2_n12_w21, 
            w22=> c2_n12_w22, 
            w23=> c2_n12_w23, 
            w24=> c2_n12_w24, 
            w25=> c2_n12_w25, 
            w26=> c2_n12_w26, 
            w27=> c2_n12_w27, 
            w28=> c2_n12_w28, 
            w29=> c2_n12_w29, 
            w30=> c2_n12_w30, 
            w31=> c2_n12_w31, 
            w32=> c2_n12_w32, 
            w33=> c2_n12_w33, 
            w34=> c2_n12_w34, 
            w35=> c2_n12_w35, 
            w36=> c2_n12_w36, 
            w37=> c2_n12_w37, 
            w38=> c2_n12_w38, 
            w39=> c2_n12_w39, 
            w40=> c2_n12_w40, 
            w41=> c2_n12_w41, 
            w42=> c2_n12_w42, 
            w43=> c2_n12_w43, 
            w44=> c2_n12_w44, 
            w45=> c2_n12_w45, 
            w46=> c2_n12_w46, 
            w47=> c2_n12_w47, 
            w48=> c2_n12_w48, 
            w49=> c2_n12_w49, 
            w50=> c2_n12_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n12_y
   );           
            
neuron_inst_13: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n13_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n13_w1, 
            w2=> c2_n13_w2, 
            w3=> c2_n13_w3, 
            w4=> c2_n13_w4, 
            w5=> c2_n13_w5, 
            w6=> c2_n13_w6, 
            w7=> c2_n13_w7, 
            w8=> c2_n13_w8, 
            w9=> c2_n13_w9, 
            w10=> c2_n13_w10, 
            w11=> c2_n13_w11, 
            w12=> c2_n13_w12, 
            w13=> c2_n13_w13, 
            w14=> c2_n13_w14, 
            w15=> c2_n13_w15, 
            w16=> c2_n13_w16, 
            w17=> c2_n13_w17, 
            w18=> c2_n13_w18, 
            w19=> c2_n13_w19, 
            w20=> c2_n13_w20, 
            w21=> c2_n13_w21, 
            w22=> c2_n13_w22, 
            w23=> c2_n13_w23, 
            w24=> c2_n13_w24, 
            w25=> c2_n13_w25, 
            w26=> c2_n13_w26, 
            w27=> c2_n13_w27, 
            w28=> c2_n13_w28, 
            w29=> c2_n13_w29, 
            w30=> c2_n13_w30, 
            w31=> c2_n13_w31, 
            w32=> c2_n13_w32, 
            w33=> c2_n13_w33, 
            w34=> c2_n13_w34, 
            w35=> c2_n13_w35, 
            w36=> c2_n13_w36, 
            w37=> c2_n13_w37, 
            w38=> c2_n13_w38, 
            w39=> c2_n13_w39, 
            w40=> c2_n13_w40, 
            w41=> c2_n13_w41, 
            w42=> c2_n13_w42, 
            w43=> c2_n13_w43, 
            w44=> c2_n13_w44, 
            w45=> c2_n13_w45, 
            w46=> c2_n13_w46, 
            w47=> c2_n13_w47, 
            w48=> c2_n13_w48, 
            w49=> c2_n13_w49, 
            w50=> c2_n13_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n13_y
   );           
            
neuron_inst_14: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n14_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n14_w1, 
            w2=> c2_n14_w2, 
            w3=> c2_n14_w3, 
            w4=> c2_n14_w4, 
            w5=> c2_n14_w5, 
            w6=> c2_n14_w6, 
            w7=> c2_n14_w7, 
            w8=> c2_n14_w8, 
            w9=> c2_n14_w9, 
            w10=> c2_n14_w10, 
            w11=> c2_n14_w11, 
            w12=> c2_n14_w12, 
            w13=> c2_n14_w13, 
            w14=> c2_n14_w14, 
            w15=> c2_n14_w15, 
            w16=> c2_n14_w16, 
            w17=> c2_n14_w17, 
            w18=> c2_n14_w18, 
            w19=> c2_n14_w19, 
            w20=> c2_n14_w20, 
            w21=> c2_n14_w21, 
            w22=> c2_n14_w22, 
            w23=> c2_n14_w23, 
            w24=> c2_n14_w24, 
            w25=> c2_n14_w25, 
            w26=> c2_n14_w26, 
            w27=> c2_n14_w27, 
            w28=> c2_n14_w28, 
            w29=> c2_n14_w29, 
            w30=> c2_n14_w30, 
            w31=> c2_n14_w31, 
            w32=> c2_n14_w32, 
            w33=> c2_n14_w33, 
            w34=> c2_n14_w34, 
            w35=> c2_n14_w35, 
            w36=> c2_n14_w36, 
            w37=> c2_n14_w37, 
            w38=> c2_n14_w38, 
            w39=> c2_n14_w39, 
            w40=> c2_n14_w40, 
            w41=> c2_n14_w41, 
            w42=> c2_n14_w42, 
            w43=> c2_n14_w43, 
            w44=> c2_n14_w44, 
            w45=> c2_n14_w45, 
            w46=> c2_n14_w46, 
            w47=> c2_n14_w47, 
            w48=> c2_n14_w48, 
            w49=> c2_n14_w49, 
            w50=> c2_n14_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n14_y
   );           
            
neuron_inst_15: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n15_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n15_w1, 
            w2=> c2_n15_w2, 
            w3=> c2_n15_w3, 
            w4=> c2_n15_w4, 
            w5=> c2_n15_w5, 
            w6=> c2_n15_w6, 
            w7=> c2_n15_w7, 
            w8=> c2_n15_w8, 
            w9=> c2_n15_w9, 
            w10=> c2_n15_w10, 
            w11=> c2_n15_w11, 
            w12=> c2_n15_w12, 
            w13=> c2_n15_w13, 
            w14=> c2_n15_w14, 
            w15=> c2_n15_w15, 
            w16=> c2_n15_w16, 
            w17=> c2_n15_w17, 
            w18=> c2_n15_w18, 
            w19=> c2_n15_w19, 
            w20=> c2_n15_w20, 
            w21=> c2_n15_w21, 
            w22=> c2_n15_w22, 
            w23=> c2_n15_w23, 
            w24=> c2_n15_w24, 
            w25=> c2_n15_w25, 
            w26=> c2_n15_w26, 
            w27=> c2_n15_w27, 
            w28=> c2_n15_w28, 
            w29=> c2_n15_w29, 
            w30=> c2_n15_w30, 
            w31=> c2_n15_w31, 
            w32=> c2_n15_w32, 
            w33=> c2_n15_w33, 
            w34=> c2_n15_w34, 
            w35=> c2_n15_w35, 
            w36=> c2_n15_w36, 
            w37=> c2_n15_w37, 
            w38=> c2_n15_w38, 
            w39=> c2_n15_w39, 
            w40=> c2_n15_w40, 
            w41=> c2_n15_w41, 
            w42=> c2_n15_w42, 
            w43=> c2_n15_w43, 
            w44=> c2_n15_w44, 
            w45=> c2_n15_w45, 
            w46=> c2_n15_w46, 
            w47=> c2_n15_w47, 
            w48=> c2_n15_w48, 
            w49=> c2_n15_w49, 
            w50=> c2_n15_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n15_y
   );           
            
neuron_inst_16: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n16_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n16_w1, 
            w2=> c2_n16_w2, 
            w3=> c2_n16_w3, 
            w4=> c2_n16_w4, 
            w5=> c2_n16_w5, 
            w6=> c2_n16_w6, 
            w7=> c2_n16_w7, 
            w8=> c2_n16_w8, 
            w9=> c2_n16_w9, 
            w10=> c2_n16_w10, 
            w11=> c2_n16_w11, 
            w12=> c2_n16_w12, 
            w13=> c2_n16_w13, 
            w14=> c2_n16_w14, 
            w15=> c2_n16_w15, 
            w16=> c2_n16_w16, 
            w17=> c2_n16_w17, 
            w18=> c2_n16_w18, 
            w19=> c2_n16_w19, 
            w20=> c2_n16_w20, 
            w21=> c2_n16_w21, 
            w22=> c2_n16_w22, 
            w23=> c2_n16_w23, 
            w24=> c2_n16_w24, 
            w25=> c2_n16_w25, 
            w26=> c2_n16_w26, 
            w27=> c2_n16_w27, 
            w28=> c2_n16_w28, 
            w29=> c2_n16_w29, 
            w30=> c2_n16_w30, 
            w31=> c2_n16_w31, 
            w32=> c2_n16_w32, 
            w33=> c2_n16_w33, 
            w34=> c2_n16_w34, 
            w35=> c2_n16_w35, 
            w36=> c2_n16_w36, 
            w37=> c2_n16_w37, 
            w38=> c2_n16_w38, 
            w39=> c2_n16_w39, 
            w40=> c2_n16_w40, 
            w41=> c2_n16_w41, 
            w42=> c2_n16_w42, 
            w43=> c2_n16_w43, 
            w44=> c2_n16_w44, 
            w45=> c2_n16_w45, 
            w46=> c2_n16_w46, 
            w47=> c2_n16_w47, 
            w48=> c2_n16_w48, 
            w49=> c2_n16_w49, 
            w50=> c2_n16_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n16_y
   );           
            
neuron_inst_17: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n17_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n17_w1, 
            w2=> c2_n17_w2, 
            w3=> c2_n17_w3, 
            w4=> c2_n17_w4, 
            w5=> c2_n17_w5, 
            w6=> c2_n17_w6, 
            w7=> c2_n17_w7, 
            w8=> c2_n17_w8, 
            w9=> c2_n17_w9, 
            w10=> c2_n17_w10, 
            w11=> c2_n17_w11, 
            w12=> c2_n17_w12, 
            w13=> c2_n17_w13, 
            w14=> c2_n17_w14, 
            w15=> c2_n17_w15, 
            w16=> c2_n17_w16, 
            w17=> c2_n17_w17, 
            w18=> c2_n17_w18, 
            w19=> c2_n17_w19, 
            w20=> c2_n17_w20, 
            w21=> c2_n17_w21, 
            w22=> c2_n17_w22, 
            w23=> c2_n17_w23, 
            w24=> c2_n17_w24, 
            w25=> c2_n17_w25, 
            w26=> c2_n17_w26, 
            w27=> c2_n17_w27, 
            w28=> c2_n17_w28, 
            w29=> c2_n17_w29, 
            w30=> c2_n17_w30, 
            w31=> c2_n17_w31, 
            w32=> c2_n17_w32, 
            w33=> c2_n17_w33, 
            w34=> c2_n17_w34, 
            w35=> c2_n17_w35, 
            w36=> c2_n17_w36, 
            w37=> c2_n17_w37, 
            w38=> c2_n17_w38, 
            w39=> c2_n17_w39, 
            w40=> c2_n17_w40, 
            w41=> c2_n17_w41, 
            w42=> c2_n17_w42, 
            w43=> c2_n17_w43, 
            w44=> c2_n17_w44, 
            w45=> c2_n17_w45, 
            w46=> c2_n17_w46, 
            w47=> c2_n17_w47, 
            w48=> c2_n17_w48, 
            w49=> c2_n17_w49, 
            w50=> c2_n17_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n17_y
   );           
            
neuron_inst_18: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n18_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n18_w1, 
            w2=> c2_n18_w2, 
            w3=> c2_n18_w3, 
            w4=> c2_n18_w4, 
            w5=> c2_n18_w5, 
            w6=> c2_n18_w6, 
            w7=> c2_n18_w7, 
            w8=> c2_n18_w8, 
            w9=> c2_n18_w9, 
            w10=> c2_n18_w10, 
            w11=> c2_n18_w11, 
            w12=> c2_n18_w12, 
            w13=> c2_n18_w13, 
            w14=> c2_n18_w14, 
            w15=> c2_n18_w15, 
            w16=> c2_n18_w16, 
            w17=> c2_n18_w17, 
            w18=> c2_n18_w18, 
            w19=> c2_n18_w19, 
            w20=> c2_n18_w20, 
            w21=> c2_n18_w21, 
            w22=> c2_n18_w22, 
            w23=> c2_n18_w23, 
            w24=> c2_n18_w24, 
            w25=> c2_n18_w25, 
            w26=> c2_n18_w26, 
            w27=> c2_n18_w27, 
            w28=> c2_n18_w28, 
            w29=> c2_n18_w29, 
            w30=> c2_n18_w30, 
            w31=> c2_n18_w31, 
            w32=> c2_n18_w32, 
            w33=> c2_n18_w33, 
            w34=> c2_n18_w34, 
            w35=> c2_n18_w35, 
            w36=> c2_n18_w36, 
            w37=> c2_n18_w37, 
            w38=> c2_n18_w38, 
            w39=> c2_n18_w39, 
            w40=> c2_n18_w40, 
            w41=> c2_n18_w41, 
            w42=> c2_n18_w42, 
            w43=> c2_n18_w43, 
            w44=> c2_n18_w44, 
            w45=> c2_n18_w45, 
            w46=> c2_n18_w46, 
            w47=> c2_n18_w47, 
            w48=> c2_n18_w48, 
            w49=> c2_n18_w49, 
            w50=> c2_n18_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n18_y
   );           
            
neuron_inst_19: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n19_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n19_w1, 
            w2=> c2_n19_w2, 
            w3=> c2_n19_w3, 
            w4=> c2_n19_w4, 
            w5=> c2_n19_w5, 
            w6=> c2_n19_w6, 
            w7=> c2_n19_w7, 
            w8=> c2_n19_w8, 
            w9=> c2_n19_w9, 
            w10=> c2_n19_w10, 
            w11=> c2_n19_w11, 
            w12=> c2_n19_w12, 
            w13=> c2_n19_w13, 
            w14=> c2_n19_w14, 
            w15=> c2_n19_w15, 
            w16=> c2_n19_w16, 
            w17=> c2_n19_w17, 
            w18=> c2_n19_w18, 
            w19=> c2_n19_w19, 
            w20=> c2_n19_w20, 
            w21=> c2_n19_w21, 
            w22=> c2_n19_w22, 
            w23=> c2_n19_w23, 
            w24=> c2_n19_w24, 
            w25=> c2_n19_w25, 
            w26=> c2_n19_w26, 
            w27=> c2_n19_w27, 
            w28=> c2_n19_w28, 
            w29=> c2_n19_w29, 
            w30=> c2_n19_w30, 
            w31=> c2_n19_w31, 
            w32=> c2_n19_w32, 
            w33=> c2_n19_w33, 
            w34=> c2_n19_w34, 
            w35=> c2_n19_w35, 
            w36=> c2_n19_w36, 
            w37=> c2_n19_w37, 
            w38=> c2_n19_w38, 
            w39=> c2_n19_w39, 
            w40=> c2_n19_w40, 
            w41=> c2_n19_w41, 
            w42=> c2_n19_w42, 
            w43=> c2_n19_w43, 
            w44=> c2_n19_w44, 
            w45=> c2_n19_w45, 
            w46=> c2_n19_w46, 
            w47=> c2_n19_w47, 
            w48=> c2_n19_w48, 
            w49=> c2_n19_w49, 
            w50=> c2_n19_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n19_y
   );           
            
neuron_inst_20: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n20_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n20_w1, 
            w2=> c2_n20_w2, 
            w3=> c2_n20_w3, 
            w4=> c2_n20_w4, 
            w5=> c2_n20_w5, 
            w6=> c2_n20_w6, 
            w7=> c2_n20_w7, 
            w8=> c2_n20_w8, 
            w9=> c2_n20_w9, 
            w10=> c2_n20_w10, 
            w11=> c2_n20_w11, 
            w12=> c2_n20_w12, 
            w13=> c2_n20_w13, 
            w14=> c2_n20_w14, 
            w15=> c2_n20_w15, 
            w16=> c2_n20_w16, 
            w17=> c2_n20_w17, 
            w18=> c2_n20_w18, 
            w19=> c2_n20_w19, 
            w20=> c2_n20_w20, 
            w21=> c2_n20_w21, 
            w22=> c2_n20_w22, 
            w23=> c2_n20_w23, 
            w24=> c2_n20_w24, 
            w25=> c2_n20_w25, 
            w26=> c2_n20_w26, 
            w27=> c2_n20_w27, 
            w28=> c2_n20_w28, 
            w29=> c2_n20_w29, 
            w30=> c2_n20_w30, 
            w31=> c2_n20_w31, 
            w32=> c2_n20_w32, 
            w33=> c2_n20_w33, 
            w34=> c2_n20_w34, 
            w35=> c2_n20_w35, 
            w36=> c2_n20_w36, 
            w37=> c2_n20_w37, 
            w38=> c2_n20_w38, 
            w39=> c2_n20_w39, 
            w40=> c2_n20_w40, 
            w41=> c2_n20_w41, 
            w42=> c2_n20_w42, 
            w43=> c2_n20_w43, 
            w44=> c2_n20_w44, 
            w45=> c2_n20_w45, 
            w46=> c2_n20_w46, 
            w47=> c2_n20_w47, 
            w48=> c2_n20_w48, 
            w49=> c2_n20_w49, 
            w50=> c2_n20_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n20_y
   );           
            
neuron_inst_21: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n21_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n21_w1, 
            w2=> c2_n21_w2, 
            w3=> c2_n21_w3, 
            w4=> c2_n21_w4, 
            w5=> c2_n21_w5, 
            w6=> c2_n21_w6, 
            w7=> c2_n21_w7, 
            w8=> c2_n21_w8, 
            w9=> c2_n21_w9, 
            w10=> c2_n21_w10, 
            w11=> c2_n21_w11, 
            w12=> c2_n21_w12, 
            w13=> c2_n21_w13, 
            w14=> c2_n21_w14, 
            w15=> c2_n21_w15, 
            w16=> c2_n21_w16, 
            w17=> c2_n21_w17, 
            w18=> c2_n21_w18, 
            w19=> c2_n21_w19, 
            w20=> c2_n21_w20, 
            w21=> c2_n21_w21, 
            w22=> c2_n21_w22, 
            w23=> c2_n21_w23, 
            w24=> c2_n21_w24, 
            w25=> c2_n21_w25, 
            w26=> c2_n21_w26, 
            w27=> c2_n21_w27, 
            w28=> c2_n21_w28, 
            w29=> c2_n21_w29, 
            w30=> c2_n21_w30, 
            w31=> c2_n21_w31, 
            w32=> c2_n21_w32, 
            w33=> c2_n21_w33, 
            w34=> c2_n21_w34, 
            w35=> c2_n21_w35, 
            w36=> c2_n21_w36, 
            w37=> c2_n21_w37, 
            w38=> c2_n21_w38, 
            w39=> c2_n21_w39, 
            w40=> c2_n21_w40, 
            w41=> c2_n21_w41, 
            w42=> c2_n21_w42, 
            w43=> c2_n21_w43, 
            w44=> c2_n21_w44, 
            w45=> c2_n21_w45, 
            w46=> c2_n21_w46, 
            w47=> c2_n21_w47, 
            w48=> c2_n21_w48, 
            w49=> c2_n21_w49, 
            w50=> c2_n21_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n21_y
   );           
            
neuron_inst_22: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n22_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n22_w1, 
            w2=> c2_n22_w2, 
            w3=> c2_n22_w3, 
            w4=> c2_n22_w4, 
            w5=> c2_n22_w5, 
            w6=> c2_n22_w6, 
            w7=> c2_n22_w7, 
            w8=> c2_n22_w8, 
            w9=> c2_n22_w9, 
            w10=> c2_n22_w10, 
            w11=> c2_n22_w11, 
            w12=> c2_n22_w12, 
            w13=> c2_n22_w13, 
            w14=> c2_n22_w14, 
            w15=> c2_n22_w15, 
            w16=> c2_n22_w16, 
            w17=> c2_n22_w17, 
            w18=> c2_n22_w18, 
            w19=> c2_n22_w19, 
            w20=> c2_n22_w20, 
            w21=> c2_n22_w21, 
            w22=> c2_n22_w22, 
            w23=> c2_n22_w23, 
            w24=> c2_n22_w24, 
            w25=> c2_n22_w25, 
            w26=> c2_n22_w26, 
            w27=> c2_n22_w27, 
            w28=> c2_n22_w28, 
            w29=> c2_n22_w29, 
            w30=> c2_n22_w30, 
            w31=> c2_n22_w31, 
            w32=> c2_n22_w32, 
            w33=> c2_n22_w33, 
            w34=> c2_n22_w34, 
            w35=> c2_n22_w35, 
            w36=> c2_n22_w36, 
            w37=> c2_n22_w37, 
            w38=> c2_n22_w38, 
            w39=> c2_n22_w39, 
            w40=> c2_n22_w40, 
            w41=> c2_n22_w41, 
            w42=> c2_n22_w42, 
            w43=> c2_n22_w43, 
            w44=> c2_n22_w44, 
            w45=> c2_n22_w45, 
            w46=> c2_n22_w46, 
            w47=> c2_n22_w47, 
            w48=> c2_n22_w48, 
            w49=> c2_n22_w49, 
            w50=> c2_n22_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n22_y
   );           
            
neuron_inst_23: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n23_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n23_w1, 
            w2=> c2_n23_w2, 
            w3=> c2_n23_w3, 
            w4=> c2_n23_w4, 
            w5=> c2_n23_w5, 
            w6=> c2_n23_w6, 
            w7=> c2_n23_w7, 
            w8=> c2_n23_w8, 
            w9=> c2_n23_w9, 
            w10=> c2_n23_w10, 
            w11=> c2_n23_w11, 
            w12=> c2_n23_w12, 
            w13=> c2_n23_w13, 
            w14=> c2_n23_w14, 
            w15=> c2_n23_w15, 
            w16=> c2_n23_w16, 
            w17=> c2_n23_w17, 
            w18=> c2_n23_w18, 
            w19=> c2_n23_w19, 
            w20=> c2_n23_w20, 
            w21=> c2_n23_w21, 
            w22=> c2_n23_w22, 
            w23=> c2_n23_w23, 
            w24=> c2_n23_w24, 
            w25=> c2_n23_w25, 
            w26=> c2_n23_w26, 
            w27=> c2_n23_w27, 
            w28=> c2_n23_w28, 
            w29=> c2_n23_w29, 
            w30=> c2_n23_w30, 
            w31=> c2_n23_w31, 
            w32=> c2_n23_w32, 
            w33=> c2_n23_w33, 
            w34=> c2_n23_w34, 
            w35=> c2_n23_w35, 
            w36=> c2_n23_w36, 
            w37=> c2_n23_w37, 
            w38=> c2_n23_w38, 
            w39=> c2_n23_w39, 
            w40=> c2_n23_w40, 
            w41=> c2_n23_w41, 
            w42=> c2_n23_w42, 
            w43=> c2_n23_w43, 
            w44=> c2_n23_w44, 
            w45=> c2_n23_w45, 
            w46=> c2_n23_w46, 
            w47=> c2_n23_w47, 
            w48=> c2_n23_w48, 
            w49=> c2_n23_w49, 
            w50=> c2_n23_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n23_y
   );           
            
neuron_inst_24: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n24_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n24_w1, 
            w2=> c2_n24_w2, 
            w3=> c2_n24_w3, 
            w4=> c2_n24_w4, 
            w5=> c2_n24_w5, 
            w6=> c2_n24_w6, 
            w7=> c2_n24_w7, 
            w8=> c2_n24_w8, 
            w9=> c2_n24_w9, 
            w10=> c2_n24_w10, 
            w11=> c2_n24_w11, 
            w12=> c2_n24_w12, 
            w13=> c2_n24_w13, 
            w14=> c2_n24_w14, 
            w15=> c2_n24_w15, 
            w16=> c2_n24_w16, 
            w17=> c2_n24_w17, 
            w18=> c2_n24_w18, 
            w19=> c2_n24_w19, 
            w20=> c2_n24_w20, 
            w21=> c2_n24_w21, 
            w22=> c2_n24_w22, 
            w23=> c2_n24_w23, 
            w24=> c2_n24_w24, 
            w25=> c2_n24_w25, 
            w26=> c2_n24_w26, 
            w27=> c2_n24_w27, 
            w28=> c2_n24_w28, 
            w29=> c2_n24_w29, 
            w30=> c2_n24_w30, 
            w31=> c2_n24_w31, 
            w32=> c2_n24_w32, 
            w33=> c2_n24_w33, 
            w34=> c2_n24_w34, 
            w35=> c2_n24_w35, 
            w36=> c2_n24_w36, 
            w37=> c2_n24_w37, 
            w38=> c2_n24_w38, 
            w39=> c2_n24_w39, 
            w40=> c2_n24_w40, 
            w41=> c2_n24_w41, 
            w42=> c2_n24_w42, 
            w43=> c2_n24_w43, 
            w44=> c2_n24_w44, 
            w45=> c2_n24_w45, 
            w46=> c2_n24_w46, 
            w47=> c2_n24_w47, 
            w48=> c2_n24_w48, 
            w49=> c2_n24_w49, 
            w50=> c2_n24_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n24_y
   );           
            
neuron_inst_25: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n25_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n25_w1, 
            w2=> c2_n25_w2, 
            w3=> c2_n25_w3, 
            w4=> c2_n25_w4, 
            w5=> c2_n25_w5, 
            w6=> c2_n25_w6, 
            w7=> c2_n25_w7, 
            w8=> c2_n25_w8, 
            w9=> c2_n25_w9, 
            w10=> c2_n25_w10, 
            w11=> c2_n25_w11, 
            w12=> c2_n25_w12, 
            w13=> c2_n25_w13, 
            w14=> c2_n25_w14, 
            w15=> c2_n25_w15, 
            w16=> c2_n25_w16, 
            w17=> c2_n25_w17, 
            w18=> c2_n25_w18, 
            w19=> c2_n25_w19, 
            w20=> c2_n25_w20, 
            w21=> c2_n25_w21, 
            w22=> c2_n25_w22, 
            w23=> c2_n25_w23, 
            w24=> c2_n25_w24, 
            w25=> c2_n25_w25, 
            w26=> c2_n25_w26, 
            w27=> c2_n25_w27, 
            w28=> c2_n25_w28, 
            w29=> c2_n25_w29, 
            w30=> c2_n25_w30, 
            w31=> c2_n25_w31, 
            w32=> c2_n25_w32, 
            w33=> c2_n25_w33, 
            w34=> c2_n25_w34, 
            w35=> c2_n25_w35, 
            w36=> c2_n25_w36, 
            w37=> c2_n25_w37, 
            w38=> c2_n25_w38, 
            w39=> c2_n25_w39, 
            w40=> c2_n25_w40, 
            w41=> c2_n25_w41, 
            w42=> c2_n25_w42, 
            w43=> c2_n25_w43, 
            w44=> c2_n25_w44, 
            w45=> c2_n25_w45, 
            w46=> c2_n25_w46, 
            w47=> c2_n25_w47, 
            w48=> c2_n25_w48, 
            w49=> c2_n25_w49, 
            w50=> c2_n25_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n25_y
   );           
            
neuron_inst_26: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n26_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n26_w1, 
            w2=> c2_n26_w2, 
            w3=> c2_n26_w3, 
            w4=> c2_n26_w4, 
            w5=> c2_n26_w5, 
            w6=> c2_n26_w6, 
            w7=> c2_n26_w7, 
            w8=> c2_n26_w8, 
            w9=> c2_n26_w9, 
            w10=> c2_n26_w10, 
            w11=> c2_n26_w11, 
            w12=> c2_n26_w12, 
            w13=> c2_n26_w13, 
            w14=> c2_n26_w14, 
            w15=> c2_n26_w15, 
            w16=> c2_n26_w16, 
            w17=> c2_n26_w17, 
            w18=> c2_n26_w18, 
            w19=> c2_n26_w19, 
            w20=> c2_n26_w20, 
            w21=> c2_n26_w21, 
            w22=> c2_n26_w22, 
            w23=> c2_n26_w23, 
            w24=> c2_n26_w24, 
            w25=> c2_n26_w25, 
            w26=> c2_n26_w26, 
            w27=> c2_n26_w27, 
            w28=> c2_n26_w28, 
            w29=> c2_n26_w29, 
            w30=> c2_n26_w30, 
            w31=> c2_n26_w31, 
            w32=> c2_n26_w32, 
            w33=> c2_n26_w33, 
            w34=> c2_n26_w34, 
            w35=> c2_n26_w35, 
            w36=> c2_n26_w36, 
            w37=> c2_n26_w37, 
            w38=> c2_n26_w38, 
            w39=> c2_n26_w39, 
            w40=> c2_n26_w40, 
            w41=> c2_n26_w41, 
            w42=> c2_n26_w42, 
            w43=> c2_n26_w43, 
            w44=> c2_n26_w44, 
            w45=> c2_n26_w45, 
            w46=> c2_n26_w46, 
            w47=> c2_n26_w47, 
            w48=> c2_n26_w48, 
            w49=> c2_n26_w49, 
            w50=> c2_n26_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n26_y
   );           
            
neuron_inst_27: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n27_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n27_w1, 
            w2=> c2_n27_w2, 
            w3=> c2_n27_w3, 
            w4=> c2_n27_w4, 
            w5=> c2_n27_w5, 
            w6=> c2_n27_w6, 
            w7=> c2_n27_w7, 
            w8=> c2_n27_w8, 
            w9=> c2_n27_w9, 
            w10=> c2_n27_w10, 
            w11=> c2_n27_w11, 
            w12=> c2_n27_w12, 
            w13=> c2_n27_w13, 
            w14=> c2_n27_w14, 
            w15=> c2_n27_w15, 
            w16=> c2_n27_w16, 
            w17=> c2_n27_w17, 
            w18=> c2_n27_w18, 
            w19=> c2_n27_w19, 
            w20=> c2_n27_w20, 
            w21=> c2_n27_w21, 
            w22=> c2_n27_w22, 
            w23=> c2_n27_w23, 
            w24=> c2_n27_w24, 
            w25=> c2_n27_w25, 
            w26=> c2_n27_w26, 
            w27=> c2_n27_w27, 
            w28=> c2_n27_w28, 
            w29=> c2_n27_w29, 
            w30=> c2_n27_w30, 
            w31=> c2_n27_w31, 
            w32=> c2_n27_w32, 
            w33=> c2_n27_w33, 
            w34=> c2_n27_w34, 
            w35=> c2_n27_w35, 
            w36=> c2_n27_w36, 
            w37=> c2_n27_w37, 
            w38=> c2_n27_w38, 
            w39=> c2_n27_w39, 
            w40=> c2_n27_w40, 
            w41=> c2_n27_w41, 
            w42=> c2_n27_w42, 
            w43=> c2_n27_w43, 
            w44=> c2_n27_w44, 
            w45=> c2_n27_w45, 
            w46=> c2_n27_w46, 
            w47=> c2_n27_w47, 
            w48=> c2_n27_w48, 
            w49=> c2_n27_w49, 
            w50=> c2_n27_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n27_y
   );           
            
neuron_inst_28: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n28_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n28_w1, 
            w2=> c2_n28_w2, 
            w3=> c2_n28_w3, 
            w4=> c2_n28_w4, 
            w5=> c2_n28_w5, 
            w6=> c2_n28_w6, 
            w7=> c2_n28_w7, 
            w8=> c2_n28_w8, 
            w9=> c2_n28_w9, 
            w10=> c2_n28_w10, 
            w11=> c2_n28_w11, 
            w12=> c2_n28_w12, 
            w13=> c2_n28_w13, 
            w14=> c2_n28_w14, 
            w15=> c2_n28_w15, 
            w16=> c2_n28_w16, 
            w17=> c2_n28_w17, 
            w18=> c2_n28_w18, 
            w19=> c2_n28_w19, 
            w20=> c2_n28_w20, 
            w21=> c2_n28_w21, 
            w22=> c2_n28_w22, 
            w23=> c2_n28_w23, 
            w24=> c2_n28_w24, 
            w25=> c2_n28_w25, 
            w26=> c2_n28_w26, 
            w27=> c2_n28_w27, 
            w28=> c2_n28_w28, 
            w29=> c2_n28_w29, 
            w30=> c2_n28_w30, 
            w31=> c2_n28_w31, 
            w32=> c2_n28_w32, 
            w33=> c2_n28_w33, 
            w34=> c2_n28_w34, 
            w35=> c2_n28_w35, 
            w36=> c2_n28_w36, 
            w37=> c2_n28_w37, 
            w38=> c2_n28_w38, 
            w39=> c2_n28_w39, 
            w40=> c2_n28_w40, 
            w41=> c2_n28_w41, 
            w42=> c2_n28_w42, 
            w43=> c2_n28_w43, 
            w44=> c2_n28_w44, 
            w45=> c2_n28_w45, 
            w46=> c2_n28_w46, 
            w47=> c2_n28_w47, 
            w48=> c2_n28_w48, 
            w49=> c2_n28_w49, 
            w50=> c2_n28_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n28_y
   );           
            
neuron_inst_29: ENTITY work.neuron_comb_ReLU_50n_8bit_unsigned_mul0_v0_add0_v0
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c2_n29_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            w1=> c2_n29_w1, 
            w2=> c2_n29_w2, 
            w3=> c2_n29_w3, 
            w4=> c2_n29_w4, 
            w5=> c2_n29_w5, 
            w6=> c2_n29_w6, 
            w7=> c2_n29_w7, 
            w8=> c2_n29_w8, 
            w9=> c2_n29_w9, 
            w10=> c2_n29_w10, 
            w11=> c2_n29_w11, 
            w12=> c2_n29_w12, 
            w13=> c2_n29_w13, 
            w14=> c2_n29_w14, 
            w15=> c2_n29_w15, 
            w16=> c2_n29_w16, 
            w17=> c2_n29_w17, 
            w18=> c2_n29_w18, 
            w19=> c2_n29_w19, 
            w20=> c2_n29_w20, 
            w21=> c2_n29_w21, 
            w22=> c2_n29_w22, 
            w23=> c2_n29_w23, 
            w24=> c2_n29_w24, 
            w25=> c2_n29_w25, 
            w26=> c2_n29_w26, 
            w27=> c2_n29_w27, 
            w28=> c2_n29_w28, 
            w29=> c2_n29_w29, 
            w30=> c2_n29_w30, 
            w31=> c2_n29_w31, 
            w32=> c2_n29_w32, 
            w33=> c2_n29_w33, 
            w34=> c2_n29_w34, 
            w35=> c2_n29_w35, 
            w36=> c2_n29_w36, 
            w37=> c2_n29_w37, 
            w38=> c2_n29_w38, 
            w39=> c2_n29_w39, 
            w40=> c2_n29_w40, 
            w41=> c2_n29_w41, 
            w42=> c2_n29_w42, 
            w43=> c2_n29_w43, 
            w44=> c2_n29_w44, 
            w45=> c2_n29_w45, 
            w46=> c2_n29_w46, 
            w47=> c2_n29_w47, 
            w48=> c2_n29_w48, 
            w49=> c2_n29_w49, 
            w50=> c2_n29_w50, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c2_n29_y
   );           
             
END ARCHITECTURE;
