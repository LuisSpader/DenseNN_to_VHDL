LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada0_Leaky_ReLU_100neuron_8bits_75n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c0_n0_bias, c0_n1_bias, c0_n2_bias, c0_n3_bias, c0_n4_bias, c0_n5_bias, c0_n6_bias, c0_n7_bias, c0_n8_bias, c0_n9_bias, c0_n10_bias, c0_n11_bias, c0_n12_bias, c0_n13_bias, c0_n14_bias, c0_n15_bias, c0_n16_bias, c0_n17_bias, c0_n18_bias, c0_n19_bias, c0_n20_bias, c0_n21_bias, c0_n22_bias, c0_n23_bias, c0_n24_bias, c0_n25_bias, c0_n26_bias, c0_n27_bias, c0_n28_bias, c0_n29_bias, c0_n30_bias, c0_n31_bias, c0_n32_bias, c0_n33_bias, c0_n34_bias, c0_n35_bias, c0_n36_bias, c0_n37_bias, c0_n38_bias, c0_n39_bias, c0_n40_bias, c0_n41_bias, c0_n42_bias, c0_n43_bias, c0_n44_bias, c0_n45_bias, c0_n46_bias, c0_n47_bias, c0_n48_bias, c0_n49_bias, c0_n50_bias, c0_n51_bias, c0_n52_bias, c0_n53_bias, c0_n54_bias, c0_n55_bias, c0_n56_bias, c0_n57_bias, c0_n58_bias, c0_n59_bias, c0_n60_bias, c0_n61_bias, c0_n62_bias, c0_n63_bias, c0_n64_bias, c0_n65_bias, c0_n66_bias, c0_n67_bias, c0_n68_bias, c0_n69_bias, c0_n70_bias, c0_n71_bias, c0_n72_bias, c0_n73_bias, c0_n74_bias, c0_n75_bias, c0_n76_bias, c0_n77_bias, c0_n78_bias, c0_n79_bias, c0_n80_bias, c0_n81_bias, c0_n82_bias, c0_n83_bias, c0_n84_bias, c0_n85_bias, c0_n86_bias, c0_n87_bias, c0_n88_bias, c0_n89_bias, c0_n90_bias, c0_n91_bias, c0_n92_bias, c0_n93_bias, c0_n94_bias, c0_n95_bias, c0_n96_bias, c0_n97_bias, c0_n98_bias, c0_n99_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, c0_n0_w1, c0_n0_w2, c0_n0_w3, c0_n0_w4, c0_n0_w5, c0_n0_w6, c0_n0_w7, c0_n0_w8, c0_n0_w9, c0_n0_w10, c0_n0_w11, c0_n0_w12, c0_n0_w13, c0_n0_w14, c0_n0_w15, c0_n0_w16, c0_n0_w17, c0_n0_w18, c0_n0_w19, c0_n0_w20, c0_n0_w21, c0_n0_w22, c0_n0_w23, c0_n0_w24, c0_n0_w25, c0_n0_w26, c0_n0_w27, c0_n0_w28, c0_n0_w29, c0_n0_w30, c0_n0_w31, c0_n0_w32, c0_n0_w33, c0_n0_w34, c0_n0_w35, c0_n0_w36, c0_n0_w37, c0_n0_w38, c0_n0_w39, c0_n0_w40, c0_n0_w41, c0_n0_w42, c0_n0_w43, c0_n0_w44, c0_n0_w45, c0_n0_w46, c0_n0_w47, c0_n0_w48, c0_n0_w49, c0_n0_w50, c0_n0_w51, c0_n0_w52, c0_n0_w53, c0_n0_w54, c0_n0_w55, c0_n0_w56, c0_n0_w57, c0_n0_w58, c0_n0_w59, c0_n0_w60, c0_n0_w61, c0_n0_w62, c0_n0_w63, c0_n0_w64, c0_n0_w65, c0_n0_w66, c0_n0_w67, c0_n0_w68, c0_n0_w69, c0_n0_w70, c0_n0_w71, c0_n0_w72, c0_n0_w73, c0_n0_w74, c0_n0_w75, c0_n1_w1, c0_n1_w2, c0_n1_w3, c0_n1_w4, c0_n1_w5, c0_n1_w6, c0_n1_w7, c0_n1_w8, c0_n1_w9, c0_n1_w10, c0_n1_w11, c0_n1_w12, c0_n1_w13, c0_n1_w14, c0_n1_w15, c0_n1_w16, c0_n1_w17, c0_n1_w18, c0_n1_w19, c0_n1_w20, c0_n1_w21, c0_n1_w22, c0_n1_w23, c0_n1_w24, c0_n1_w25, c0_n1_w26, c0_n1_w27, c0_n1_w28, c0_n1_w29, c0_n1_w30, c0_n1_w31, c0_n1_w32, c0_n1_w33, c0_n1_w34, c0_n1_w35, c0_n1_w36, c0_n1_w37, c0_n1_w38, c0_n1_w39, c0_n1_w40, c0_n1_w41, c0_n1_w42, c0_n1_w43, c0_n1_w44, c0_n1_w45, c0_n1_w46, c0_n1_w47, c0_n1_w48, c0_n1_w49, c0_n1_w50, c0_n1_w51, c0_n1_w52, c0_n1_w53, c0_n1_w54, c0_n1_w55, c0_n1_w56, c0_n1_w57, c0_n1_w58, c0_n1_w59, c0_n1_w60, c0_n1_w61, c0_n1_w62, c0_n1_w63, c0_n1_w64, c0_n1_w65, c0_n1_w66, c0_n1_w67, c0_n1_w68, c0_n1_w69, c0_n1_w70, c0_n1_w71, c0_n1_w72, c0_n1_w73, c0_n1_w74, c0_n1_w75, c0_n2_w1, c0_n2_w2, c0_n2_w3, c0_n2_w4, c0_n2_w5, c0_n2_w6, c0_n2_w7, c0_n2_w8, c0_n2_w9, c0_n2_w10, c0_n2_w11, c0_n2_w12, c0_n2_w13, c0_n2_w14, c0_n2_w15, c0_n2_w16, c0_n2_w17, c0_n2_w18, c0_n2_w19, c0_n2_w20, c0_n2_w21, c0_n2_w22, c0_n2_w23, c0_n2_w24, c0_n2_w25, c0_n2_w26, c0_n2_w27, c0_n2_w28, c0_n2_w29, c0_n2_w30, c0_n2_w31, c0_n2_w32, c0_n2_w33, c0_n2_w34, c0_n2_w35, c0_n2_w36, c0_n2_w37, c0_n2_w38, c0_n2_w39, c0_n2_w40, c0_n2_w41, c0_n2_w42, c0_n2_w43, c0_n2_w44, c0_n2_w45, c0_n2_w46, c0_n2_w47, c0_n2_w48, c0_n2_w49, c0_n2_w50, c0_n2_w51, c0_n2_w52, c0_n2_w53, c0_n2_w54, c0_n2_w55, c0_n2_w56, c0_n2_w57, c0_n2_w58, c0_n2_w59, c0_n2_w60, c0_n2_w61, c0_n2_w62, c0_n2_w63, c0_n2_w64, c0_n2_w65, c0_n2_w66, c0_n2_w67, c0_n2_w68, c0_n2_w69, c0_n2_w70, c0_n2_w71, c0_n2_w72, c0_n2_w73, c0_n2_w74, c0_n2_w75, c0_n3_w1, c0_n3_w2, c0_n3_w3, c0_n3_w4, c0_n3_w5, c0_n3_w6, c0_n3_w7, c0_n3_w8, c0_n3_w9, c0_n3_w10, c0_n3_w11, c0_n3_w12, c0_n3_w13, c0_n3_w14, c0_n3_w15, c0_n3_w16, c0_n3_w17, c0_n3_w18, c0_n3_w19, c0_n3_w20, c0_n3_w21, c0_n3_w22, c0_n3_w23, c0_n3_w24, c0_n3_w25, c0_n3_w26, c0_n3_w27, c0_n3_w28, c0_n3_w29, c0_n3_w30, c0_n3_w31, c0_n3_w32, c0_n3_w33, c0_n3_w34, c0_n3_w35, c0_n3_w36, c0_n3_w37, c0_n3_w38, c0_n3_w39, c0_n3_w40, c0_n3_w41, c0_n3_w42, c0_n3_w43, c0_n3_w44, c0_n3_w45, c0_n3_w46, c0_n3_w47, c0_n3_w48, c0_n3_w49, c0_n3_w50, c0_n3_w51, c0_n3_w52, c0_n3_w53, c0_n3_w54, c0_n3_w55, c0_n3_w56, c0_n3_w57, c0_n3_w58, c0_n3_w59, c0_n3_w60, c0_n3_w61, c0_n3_w62, c0_n3_w63, c0_n3_w64, c0_n3_w65, c0_n3_w66, c0_n3_w67, c0_n3_w68, c0_n3_w69, c0_n3_w70, c0_n3_w71, c0_n3_w72, c0_n3_w73, c0_n3_w74, c0_n3_w75, c0_n4_w1, c0_n4_w2, c0_n4_w3, c0_n4_w4, c0_n4_w5, c0_n4_w6, c0_n4_w7, c0_n4_w8, c0_n4_w9, c0_n4_w10, c0_n4_w11, c0_n4_w12, c0_n4_w13, c0_n4_w14, c0_n4_w15, c0_n4_w16, c0_n4_w17, c0_n4_w18, c0_n4_w19, c0_n4_w20, c0_n4_w21, c0_n4_w22, c0_n4_w23, c0_n4_w24, c0_n4_w25, c0_n4_w26, c0_n4_w27, c0_n4_w28, c0_n4_w29, c0_n4_w30, c0_n4_w31, c0_n4_w32, c0_n4_w33, c0_n4_w34, c0_n4_w35, c0_n4_w36, c0_n4_w37, c0_n4_w38, c0_n4_w39, c0_n4_w40, c0_n4_w41, c0_n4_w42, c0_n4_w43, c0_n4_w44, c0_n4_w45, c0_n4_w46, c0_n4_w47, c0_n4_w48, c0_n4_w49, c0_n4_w50, c0_n4_w51, c0_n4_w52, c0_n4_w53, c0_n4_w54, c0_n4_w55, c0_n4_w56, c0_n4_w57, c0_n4_w58, c0_n4_w59, c0_n4_w60, c0_n4_w61, c0_n4_w62, c0_n4_w63, c0_n4_w64, c0_n4_w65, c0_n4_w66, c0_n4_w67, c0_n4_w68, c0_n4_w69, c0_n4_w70, c0_n4_w71, c0_n4_w72, c0_n4_w73, c0_n4_w74, c0_n4_w75, c0_n5_w1, c0_n5_w2, c0_n5_w3, c0_n5_w4, c0_n5_w5, c0_n5_w6, c0_n5_w7, c0_n5_w8, c0_n5_w9, c0_n5_w10, c0_n5_w11, c0_n5_w12, c0_n5_w13, c0_n5_w14, c0_n5_w15, c0_n5_w16, c0_n5_w17, c0_n5_w18, c0_n5_w19, c0_n5_w20, c0_n5_w21, c0_n5_w22, c0_n5_w23, c0_n5_w24, c0_n5_w25, c0_n5_w26, c0_n5_w27, c0_n5_w28, c0_n5_w29, c0_n5_w30, c0_n5_w31, c0_n5_w32, c0_n5_w33, c0_n5_w34, c0_n5_w35, c0_n5_w36, c0_n5_w37, c0_n5_w38, c0_n5_w39, c0_n5_w40, c0_n5_w41, c0_n5_w42, c0_n5_w43, c0_n5_w44, c0_n5_w45, c0_n5_w46, c0_n5_w47, c0_n5_w48, c0_n5_w49, c0_n5_w50, c0_n5_w51, c0_n5_w52, c0_n5_w53, c0_n5_w54, c0_n5_w55, c0_n5_w56, c0_n5_w57, c0_n5_w58, c0_n5_w59, c0_n5_w60, c0_n5_w61, c0_n5_w62, c0_n5_w63, c0_n5_w64, c0_n5_w65, c0_n5_w66, c0_n5_w67, c0_n5_w68, c0_n5_w69, c0_n5_w70, c0_n5_w71, c0_n5_w72, c0_n5_w73, c0_n5_w74, c0_n5_w75, c0_n6_w1, c0_n6_w2, c0_n6_w3, c0_n6_w4, c0_n6_w5, c0_n6_w6, c0_n6_w7, c0_n6_w8, c0_n6_w9, c0_n6_w10, c0_n6_w11, c0_n6_w12, c0_n6_w13, c0_n6_w14, c0_n6_w15, c0_n6_w16, c0_n6_w17, c0_n6_w18, c0_n6_w19, c0_n6_w20, c0_n6_w21, c0_n6_w22, c0_n6_w23, c0_n6_w24, c0_n6_w25, c0_n6_w26, c0_n6_w27, c0_n6_w28, c0_n6_w29, c0_n6_w30, c0_n6_w31, c0_n6_w32, c0_n6_w33, c0_n6_w34, c0_n6_w35, c0_n6_w36, c0_n6_w37, c0_n6_w38, c0_n6_w39, c0_n6_w40, c0_n6_w41, c0_n6_w42, c0_n6_w43, c0_n6_w44, c0_n6_w45, c0_n6_w46, c0_n6_w47, c0_n6_w48, c0_n6_w49, c0_n6_w50, c0_n6_w51, c0_n6_w52, c0_n6_w53, c0_n6_w54, c0_n6_w55, c0_n6_w56, c0_n6_w57, c0_n6_w58, c0_n6_w59, c0_n6_w60, c0_n6_w61, c0_n6_w62, c0_n6_w63, c0_n6_w64, c0_n6_w65, c0_n6_w66, c0_n6_w67, c0_n6_w68, c0_n6_w69, c0_n6_w70, c0_n6_w71, c0_n6_w72, c0_n6_w73, c0_n6_w74, c0_n6_w75, c0_n7_w1, c0_n7_w2, c0_n7_w3, c0_n7_w4, c0_n7_w5, c0_n7_w6, c0_n7_w7, c0_n7_w8, c0_n7_w9, c0_n7_w10, c0_n7_w11, c0_n7_w12, c0_n7_w13, c0_n7_w14, c0_n7_w15, c0_n7_w16, c0_n7_w17, c0_n7_w18, c0_n7_w19, c0_n7_w20, c0_n7_w21, c0_n7_w22, c0_n7_w23, c0_n7_w24, c0_n7_w25, c0_n7_w26, c0_n7_w27, c0_n7_w28, c0_n7_w29, c0_n7_w30, c0_n7_w31, c0_n7_w32, c0_n7_w33, c0_n7_w34, c0_n7_w35, c0_n7_w36, c0_n7_w37, c0_n7_w38, c0_n7_w39, c0_n7_w40, c0_n7_w41, c0_n7_w42, c0_n7_w43, c0_n7_w44, c0_n7_w45, c0_n7_w46, c0_n7_w47, c0_n7_w48, c0_n7_w49, c0_n7_w50, c0_n7_w51, c0_n7_w52, c0_n7_w53, c0_n7_w54, c0_n7_w55, c0_n7_w56, c0_n7_w57, c0_n7_w58, c0_n7_w59, c0_n7_w60, c0_n7_w61, c0_n7_w62, c0_n7_w63, c0_n7_w64, c0_n7_w65, c0_n7_w66, c0_n7_w67, c0_n7_w68, c0_n7_w69, c0_n7_w70, c0_n7_w71, c0_n7_w72, c0_n7_w73, c0_n7_w74, c0_n7_w75, c0_n8_w1, c0_n8_w2, c0_n8_w3, c0_n8_w4, c0_n8_w5, c0_n8_w6, c0_n8_w7, c0_n8_w8, c0_n8_w9, c0_n8_w10, c0_n8_w11, c0_n8_w12, c0_n8_w13, c0_n8_w14, c0_n8_w15, c0_n8_w16, c0_n8_w17, c0_n8_w18, c0_n8_w19, c0_n8_w20, c0_n8_w21, c0_n8_w22, c0_n8_w23, c0_n8_w24, c0_n8_w25, c0_n8_w26, c0_n8_w27, c0_n8_w28, c0_n8_w29, c0_n8_w30, c0_n8_w31, c0_n8_w32, c0_n8_w33, c0_n8_w34, c0_n8_w35, c0_n8_w36, c0_n8_w37, c0_n8_w38, c0_n8_w39, c0_n8_w40, c0_n8_w41, c0_n8_w42, c0_n8_w43, c0_n8_w44, c0_n8_w45, c0_n8_w46, c0_n8_w47, c0_n8_w48, c0_n8_w49, c0_n8_w50, c0_n8_w51, c0_n8_w52, c0_n8_w53, c0_n8_w54, c0_n8_w55, c0_n8_w56, c0_n8_w57, c0_n8_w58, c0_n8_w59, c0_n8_w60, c0_n8_w61, c0_n8_w62, c0_n8_w63, c0_n8_w64, c0_n8_w65, c0_n8_w66, c0_n8_w67, c0_n8_w68, c0_n8_w69, c0_n8_w70, c0_n8_w71, c0_n8_w72, c0_n8_w73, c0_n8_w74, c0_n8_w75, c0_n9_w1, c0_n9_w2, c0_n9_w3, c0_n9_w4, c0_n9_w5, c0_n9_w6, c0_n9_w7, c0_n9_w8, c0_n9_w9, c0_n9_w10, c0_n9_w11, c0_n9_w12, c0_n9_w13, c0_n9_w14, c0_n9_w15, c0_n9_w16, c0_n9_w17, c0_n9_w18, c0_n9_w19, c0_n9_w20, c0_n9_w21, c0_n9_w22, c0_n9_w23, c0_n9_w24, c0_n9_w25, c0_n9_w26, c0_n9_w27, c0_n9_w28, c0_n9_w29, c0_n9_w30, c0_n9_w31, c0_n9_w32, c0_n9_w33, c0_n9_w34, c0_n9_w35, c0_n9_w36, c0_n9_w37, c0_n9_w38, c0_n9_w39, c0_n9_w40, c0_n9_w41, c0_n9_w42, c0_n9_w43, c0_n9_w44, c0_n9_w45, c0_n9_w46, c0_n9_w47, c0_n9_w48, c0_n9_w49, c0_n9_w50, c0_n9_w51, c0_n9_w52, c0_n9_w53, c0_n9_w54, c0_n9_w55, c0_n9_w56, c0_n9_w57, c0_n9_w58, c0_n9_w59, c0_n9_w60, c0_n9_w61, c0_n9_w62, c0_n9_w63, c0_n9_w64, c0_n9_w65, c0_n9_w66, c0_n9_w67, c0_n9_w68, c0_n9_w69, c0_n9_w70, c0_n9_w71, c0_n9_w72, c0_n9_w73, c0_n9_w74, c0_n9_w75, c0_n10_w1, c0_n10_w2, c0_n10_w3, c0_n10_w4, c0_n10_w5, c0_n10_w6, c0_n10_w7, c0_n10_w8, c0_n10_w9, c0_n10_w10, c0_n10_w11, c0_n10_w12, c0_n10_w13, c0_n10_w14, c0_n10_w15, c0_n10_w16, c0_n10_w17, c0_n10_w18, c0_n10_w19, c0_n10_w20, c0_n10_w21, c0_n10_w22, c0_n10_w23, c0_n10_w24, c0_n10_w25, c0_n10_w26, c0_n10_w27, c0_n10_w28, c0_n10_w29, c0_n10_w30, c0_n10_w31, c0_n10_w32, c0_n10_w33, c0_n10_w34, c0_n10_w35, c0_n10_w36, c0_n10_w37, c0_n10_w38, c0_n10_w39, c0_n10_w40, c0_n10_w41, c0_n10_w42, c0_n10_w43, c0_n10_w44, c0_n10_w45, c0_n10_w46, c0_n10_w47, c0_n10_w48, c0_n10_w49, c0_n10_w50, c0_n10_w51, c0_n10_w52, c0_n10_w53, c0_n10_w54, c0_n10_w55, c0_n10_w56, c0_n10_w57, c0_n10_w58, c0_n10_w59, c0_n10_w60, c0_n10_w61, c0_n10_w62, c0_n10_w63, c0_n10_w64, c0_n10_w65, c0_n10_w66, c0_n10_w67, c0_n10_w68, c0_n10_w69, c0_n10_w70, c0_n10_w71, c0_n10_w72, c0_n10_w73, c0_n10_w74, c0_n10_w75, c0_n11_w1, c0_n11_w2, c0_n11_w3, c0_n11_w4, c0_n11_w5, c0_n11_w6, c0_n11_w7, c0_n11_w8, c0_n11_w9, c0_n11_w10, c0_n11_w11, c0_n11_w12, c0_n11_w13, c0_n11_w14, c0_n11_w15, c0_n11_w16, c0_n11_w17, c0_n11_w18, c0_n11_w19, c0_n11_w20, c0_n11_w21, c0_n11_w22, c0_n11_w23, c0_n11_w24, c0_n11_w25, c0_n11_w26, c0_n11_w27, c0_n11_w28, c0_n11_w29, c0_n11_w30, c0_n11_w31, c0_n11_w32, c0_n11_w33, c0_n11_w34, c0_n11_w35, c0_n11_w36, c0_n11_w37, c0_n11_w38, c0_n11_w39, c0_n11_w40, c0_n11_w41, c0_n11_w42, c0_n11_w43, c0_n11_w44, c0_n11_w45, c0_n11_w46, c0_n11_w47, c0_n11_w48, c0_n11_w49, c0_n11_w50, c0_n11_w51, c0_n11_w52, c0_n11_w53, c0_n11_w54, c0_n11_w55, c0_n11_w56, c0_n11_w57, c0_n11_w58, c0_n11_w59, c0_n11_w60, c0_n11_w61, c0_n11_w62, c0_n11_w63, c0_n11_w64, c0_n11_w65, c0_n11_w66, c0_n11_w67, c0_n11_w68, c0_n11_w69, c0_n11_w70, c0_n11_w71, c0_n11_w72, c0_n11_w73, c0_n11_w74, c0_n11_w75, c0_n12_w1, c0_n12_w2, c0_n12_w3, c0_n12_w4, c0_n12_w5, c0_n12_w6, c0_n12_w7, c0_n12_w8, c0_n12_w9, c0_n12_w10, c0_n12_w11, c0_n12_w12, c0_n12_w13, c0_n12_w14, c0_n12_w15, c0_n12_w16, c0_n12_w17, c0_n12_w18, c0_n12_w19, c0_n12_w20, c0_n12_w21, c0_n12_w22, c0_n12_w23, c0_n12_w24, c0_n12_w25, c0_n12_w26, c0_n12_w27, c0_n12_w28, c0_n12_w29, c0_n12_w30, c0_n12_w31, c0_n12_w32, c0_n12_w33, c0_n12_w34, c0_n12_w35, c0_n12_w36, c0_n12_w37, c0_n12_w38, c0_n12_w39, c0_n12_w40, c0_n12_w41, c0_n12_w42, c0_n12_w43, c0_n12_w44, c0_n12_w45, c0_n12_w46, c0_n12_w47, c0_n12_w48, c0_n12_w49, c0_n12_w50, c0_n12_w51, c0_n12_w52, c0_n12_w53, c0_n12_w54, c0_n12_w55, c0_n12_w56, c0_n12_w57, c0_n12_w58, c0_n12_w59, c0_n12_w60, c0_n12_w61, c0_n12_w62, c0_n12_w63, c0_n12_w64, c0_n12_w65, c0_n12_w66, c0_n12_w67, c0_n12_w68, c0_n12_w69, c0_n12_w70, c0_n12_w71, c0_n12_w72, c0_n12_w73, c0_n12_w74, c0_n12_w75, c0_n13_w1, c0_n13_w2, c0_n13_w3, c0_n13_w4, c0_n13_w5, c0_n13_w6, c0_n13_w7, c0_n13_w8, c0_n13_w9, c0_n13_w10, c0_n13_w11, c0_n13_w12, c0_n13_w13, c0_n13_w14, c0_n13_w15, c0_n13_w16, c0_n13_w17, c0_n13_w18, c0_n13_w19, c0_n13_w20, c0_n13_w21, c0_n13_w22, c0_n13_w23, c0_n13_w24, c0_n13_w25, c0_n13_w26, c0_n13_w27, c0_n13_w28, c0_n13_w29, c0_n13_w30, c0_n13_w31, c0_n13_w32, c0_n13_w33, c0_n13_w34, c0_n13_w35, c0_n13_w36, c0_n13_w37, c0_n13_w38, c0_n13_w39, c0_n13_w40, c0_n13_w41, c0_n13_w42, c0_n13_w43, c0_n13_w44, c0_n13_w45, c0_n13_w46, c0_n13_w47, c0_n13_w48, c0_n13_w49, c0_n13_w50, c0_n13_w51, c0_n13_w52, c0_n13_w53, c0_n13_w54, c0_n13_w55, c0_n13_w56, c0_n13_w57, c0_n13_w58, c0_n13_w59, c0_n13_w60, c0_n13_w61, c0_n13_w62, c0_n13_w63, c0_n13_w64, c0_n13_w65, c0_n13_w66, c0_n13_w67, c0_n13_w68, c0_n13_w69, c0_n13_w70, c0_n13_w71, c0_n13_w72, c0_n13_w73, c0_n13_w74, c0_n13_w75, c0_n14_w1, c0_n14_w2, c0_n14_w3, c0_n14_w4, c0_n14_w5, c0_n14_w6, c0_n14_w7, c0_n14_w8, c0_n14_w9, c0_n14_w10, c0_n14_w11, c0_n14_w12, c0_n14_w13, c0_n14_w14, c0_n14_w15, c0_n14_w16, c0_n14_w17, c0_n14_w18, c0_n14_w19, c0_n14_w20, c0_n14_w21, c0_n14_w22, c0_n14_w23, c0_n14_w24, c0_n14_w25, c0_n14_w26, c0_n14_w27, c0_n14_w28, c0_n14_w29, c0_n14_w30, c0_n14_w31, c0_n14_w32, c0_n14_w33, c0_n14_w34, c0_n14_w35, c0_n14_w36, c0_n14_w37, c0_n14_w38, c0_n14_w39, c0_n14_w40, c0_n14_w41, c0_n14_w42, c0_n14_w43, c0_n14_w44, c0_n14_w45, c0_n14_w46, c0_n14_w47, c0_n14_w48, c0_n14_w49, c0_n14_w50, c0_n14_w51, c0_n14_w52, c0_n14_w53, c0_n14_w54, c0_n14_w55, c0_n14_w56, c0_n14_w57, c0_n14_w58, c0_n14_w59, c0_n14_w60, c0_n14_w61, c0_n14_w62, c0_n14_w63, c0_n14_w64, c0_n14_w65, c0_n14_w66, c0_n14_w67, c0_n14_w68, c0_n14_w69, c0_n14_w70, c0_n14_w71, c0_n14_w72, c0_n14_w73, c0_n14_w74, c0_n14_w75, c0_n15_w1, c0_n15_w2, c0_n15_w3, c0_n15_w4, c0_n15_w5, c0_n15_w6, c0_n15_w7, c0_n15_w8, c0_n15_w9, c0_n15_w10, c0_n15_w11, c0_n15_w12, c0_n15_w13, c0_n15_w14, c0_n15_w15, c0_n15_w16, c0_n15_w17, c0_n15_w18, c0_n15_w19, c0_n15_w20, c0_n15_w21, c0_n15_w22, c0_n15_w23, c0_n15_w24, c0_n15_w25, c0_n15_w26, c0_n15_w27, c0_n15_w28, c0_n15_w29, c0_n15_w30, c0_n15_w31, c0_n15_w32, c0_n15_w33, c0_n15_w34, c0_n15_w35, c0_n15_w36, c0_n15_w37, c0_n15_w38, c0_n15_w39, c0_n15_w40, c0_n15_w41, c0_n15_w42, c0_n15_w43, c0_n15_w44, c0_n15_w45, c0_n15_w46, c0_n15_w47, c0_n15_w48, c0_n15_w49, c0_n15_w50, c0_n15_w51, c0_n15_w52, c0_n15_w53, c0_n15_w54, c0_n15_w55, c0_n15_w56, c0_n15_w57, c0_n15_w58, c0_n15_w59, c0_n15_w60, c0_n15_w61, c0_n15_w62, c0_n15_w63, c0_n15_w64, c0_n15_w65, c0_n15_w66, c0_n15_w67, c0_n15_w68, c0_n15_w69, c0_n15_w70, c0_n15_w71, c0_n15_w72, c0_n15_w73, c0_n15_w74, c0_n15_w75, c0_n16_w1, c0_n16_w2, c0_n16_w3, c0_n16_w4, c0_n16_w5, c0_n16_w6, c0_n16_w7, c0_n16_w8, c0_n16_w9, c0_n16_w10, c0_n16_w11, c0_n16_w12, c0_n16_w13, c0_n16_w14, c0_n16_w15, c0_n16_w16, c0_n16_w17, c0_n16_w18, c0_n16_w19, c0_n16_w20, c0_n16_w21, c0_n16_w22, c0_n16_w23, c0_n16_w24, c0_n16_w25, c0_n16_w26, c0_n16_w27, c0_n16_w28, c0_n16_w29, c0_n16_w30, c0_n16_w31, c0_n16_w32, c0_n16_w33, c0_n16_w34, c0_n16_w35, c0_n16_w36, c0_n16_w37, c0_n16_w38, c0_n16_w39, c0_n16_w40, c0_n16_w41, c0_n16_w42, c0_n16_w43, c0_n16_w44, c0_n16_w45, c0_n16_w46, c0_n16_w47, c0_n16_w48, c0_n16_w49, c0_n16_w50, c0_n16_w51, c0_n16_w52, c0_n16_w53, c0_n16_w54, c0_n16_w55, c0_n16_w56, c0_n16_w57, c0_n16_w58, c0_n16_w59, c0_n16_w60, c0_n16_w61, c0_n16_w62, c0_n16_w63, c0_n16_w64, c0_n16_w65, c0_n16_w66, c0_n16_w67, c0_n16_w68, c0_n16_w69, c0_n16_w70, c0_n16_w71, c0_n16_w72, c0_n16_w73, c0_n16_w74, c0_n16_w75, c0_n17_w1, c0_n17_w2, c0_n17_w3, c0_n17_w4, c0_n17_w5, c0_n17_w6, c0_n17_w7, c0_n17_w8, c0_n17_w9, c0_n17_w10, c0_n17_w11, c0_n17_w12, c0_n17_w13, c0_n17_w14, c0_n17_w15, c0_n17_w16, c0_n17_w17, c0_n17_w18, c0_n17_w19, c0_n17_w20, c0_n17_w21, c0_n17_w22, c0_n17_w23, c0_n17_w24, c0_n17_w25, c0_n17_w26, c0_n17_w27, c0_n17_w28, c0_n17_w29, c0_n17_w30, c0_n17_w31, c0_n17_w32, c0_n17_w33, c0_n17_w34, c0_n17_w35, c0_n17_w36, c0_n17_w37, c0_n17_w38, c0_n17_w39, c0_n17_w40, c0_n17_w41, c0_n17_w42, c0_n17_w43, c0_n17_w44, c0_n17_w45, c0_n17_w46, c0_n17_w47, c0_n17_w48, c0_n17_w49, c0_n17_w50, c0_n17_w51, c0_n17_w52, c0_n17_w53, c0_n17_w54, c0_n17_w55, c0_n17_w56, c0_n17_w57, c0_n17_w58, c0_n17_w59, c0_n17_w60, c0_n17_w61, c0_n17_w62, c0_n17_w63, c0_n17_w64, c0_n17_w65, c0_n17_w66, c0_n17_w67, c0_n17_w68, c0_n17_w69, c0_n17_w70, c0_n17_w71, c0_n17_w72, c0_n17_w73, c0_n17_w74, c0_n17_w75, c0_n18_w1, c0_n18_w2, c0_n18_w3, c0_n18_w4, c0_n18_w5, c0_n18_w6, c0_n18_w7, c0_n18_w8, c0_n18_w9, c0_n18_w10, c0_n18_w11, c0_n18_w12, c0_n18_w13, c0_n18_w14, c0_n18_w15, c0_n18_w16, c0_n18_w17, c0_n18_w18, c0_n18_w19, c0_n18_w20, c0_n18_w21, c0_n18_w22, c0_n18_w23, c0_n18_w24, c0_n18_w25, c0_n18_w26, c0_n18_w27, c0_n18_w28, c0_n18_w29, c0_n18_w30, c0_n18_w31, c0_n18_w32, c0_n18_w33, c0_n18_w34, c0_n18_w35, c0_n18_w36, c0_n18_w37, c0_n18_w38, c0_n18_w39, c0_n18_w40, c0_n18_w41, c0_n18_w42, c0_n18_w43, c0_n18_w44, c0_n18_w45, c0_n18_w46, c0_n18_w47, c0_n18_w48, c0_n18_w49, c0_n18_w50, c0_n18_w51, c0_n18_w52, c0_n18_w53, c0_n18_w54, c0_n18_w55, c0_n18_w56, c0_n18_w57, c0_n18_w58, c0_n18_w59, c0_n18_w60, c0_n18_w61, c0_n18_w62, c0_n18_w63, c0_n18_w64, c0_n18_w65, c0_n18_w66, c0_n18_w67, c0_n18_w68, c0_n18_w69, c0_n18_w70, c0_n18_w71, c0_n18_w72, c0_n18_w73, c0_n18_w74, c0_n18_w75, c0_n19_w1, c0_n19_w2, c0_n19_w3, c0_n19_w4, c0_n19_w5, c0_n19_w6, c0_n19_w7, c0_n19_w8, c0_n19_w9, c0_n19_w10, c0_n19_w11, c0_n19_w12, c0_n19_w13, c0_n19_w14, c0_n19_w15, c0_n19_w16, c0_n19_w17, c0_n19_w18, c0_n19_w19, c0_n19_w20, c0_n19_w21, c0_n19_w22, c0_n19_w23, c0_n19_w24, c0_n19_w25, c0_n19_w26, c0_n19_w27, c0_n19_w28, c0_n19_w29, c0_n19_w30, c0_n19_w31, c0_n19_w32, c0_n19_w33, c0_n19_w34, c0_n19_w35, c0_n19_w36, c0_n19_w37, c0_n19_w38, c0_n19_w39, c0_n19_w40, c0_n19_w41, c0_n19_w42, c0_n19_w43, c0_n19_w44, c0_n19_w45, c0_n19_w46, c0_n19_w47, c0_n19_w48, c0_n19_w49, c0_n19_w50, c0_n19_w51, c0_n19_w52, c0_n19_w53, c0_n19_w54, c0_n19_w55, c0_n19_w56, c0_n19_w57, c0_n19_w58, c0_n19_w59, c0_n19_w60, c0_n19_w61, c0_n19_w62, c0_n19_w63, c0_n19_w64, c0_n19_w65, c0_n19_w66, c0_n19_w67, c0_n19_w68, c0_n19_w69, c0_n19_w70, c0_n19_w71, c0_n19_w72, c0_n19_w73, c0_n19_w74, c0_n19_w75, c0_n20_w1, c0_n20_w2, c0_n20_w3, c0_n20_w4, c0_n20_w5, c0_n20_w6, c0_n20_w7, c0_n20_w8, c0_n20_w9, c0_n20_w10, c0_n20_w11, c0_n20_w12, c0_n20_w13, c0_n20_w14, c0_n20_w15, c0_n20_w16, c0_n20_w17, c0_n20_w18, c0_n20_w19, c0_n20_w20, c0_n20_w21, c0_n20_w22, c0_n20_w23, c0_n20_w24, c0_n20_w25, c0_n20_w26, c0_n20_w27, c0_n20_w28, c0_n20_w29, c0_n20_w30, c0_n20_w31, c0_n20_w32, c0_n20_w33, c0_n20_w34, c0_n20_w35, c0_n20_w36, c0_n20_w37, c0_n20_w38, c0_n20_w39, c0_n20_w40, c0_n20_w41, c0_n20_w42, c0_n20_w43, c0_n20_w44, c0_n20_w45, c0_n20_w46, c0_n20_w47, c0_n20_w48, c0_n20_w49, c0_n20_w50, c0_n20_w51, c0_n20_w52, c0_n20_w53, c0_n20_w54, c0_n20_w55, c0_n20_w56, c0_n20_w57, c0_n20_w58, c0_n20_w59, c0_n20_w60, c0_n20_w61, c0_n20_w62, c0_n20_w63, c0_n20_w64, c0_n20_w65, c0_n20_w66, c0_n20_w67, c0_n20_w68, c0_n20_w69, c0_n20_w70, c0_n20_w71, c0_n20_w72, c0_n20_w73, c0_n20_w74, c0_n20_w75, c0_n21_w1, c0_n21_w2, c0_n21_w3, c0_n21_w4, c0_n21_w5, c0_n21_w6, c0_n21_w7, c0_n21_w8, c0_n21_w9, c0_n21_w10, c0_n21_w11, c0_n21_w12, c0_n21_w13, c0_n21_w14, c0_n21_w15, c0_n21_w16, c0_n21_w17, c0_n21_w18, c0_n21_w19, c0_n21_w20, c0_n21_w21, c0_n21_w22, c0_n21_w23, c0_n21_w24, c0_n21_w25, c0_n21_w26, c0_n21_w27, c0_n21_w28, c0_n21_w29, c0_n21_w30, c0_n21_w31, c0_n21_w32, c0_n21_w33, c0_n21_w34, c0_n21_w35, c0_n21_w36, c0_n21_w37, c0_n21_w38, c0_n21_w39, c0_n21_w40, c0_n21_w41, c0_n21_w42, c0_n21_w43, c0_n21_w44, c0_n21_w45, c0_n21_w46, c0_n21_w47, c0_n21_w48, c0_n21_w49, c0_n21_w50, c0_n21_w51, c0_n21_w52, c0_n21_w53, c0_n21_w54, c0_n21_w55, c0_n21_w56, c0_n21_w57, c0_n21_w58, c0_n21_w59, c0_n21_w60, c0_n21_w61, c0_n21_w62, c0_n21_w63, c0_n21_w64, c0_n21_w65, c0_n21_w66, c0_n21_w67, c0_n21_w68, c0_n21_w69, c0_n21_w70, c0_n21_w71, c0_n21_w72, c0_n21_w73, c0_n21_w74, c0_n21_w75, c0_n22_w1, c0_n22_w2, c0_n22_w3, c0_n22_w4, c0_n22_w5, c0_n22_w6, c0_n22_w7, c0_n22_w8, c0_n22_w9, c0_n22_w10, c0_n22_w11, c0_n22_w12, c0_n22_w13, c0_n22_w14, c0_n22_w15, c0_n22_w16, c0_n22_w17, c0_n22_w18, c0_n22_w19, c0_n22_w20, c0_n22_w21, c0_n22_w22, c0_n22_w23, c0_n22_w24, c0_n22_w25, c0_n22_w26, c0_n22_w27, c0_n22_w28, c0_n22_w29, c0_n22_w30, c0_n22_w31, c0_n22_w32, c0_n22_w33, c0_n22_w34, c0_n22_w35, c0_n22_w36, c0_n22_w37, c0_n22_w38, c0_n22_w39, c0_n22_w40, c0_n22_w41, c0_n22_w42, c0_n22_w43, c0_n22_w44, c0_n22_w45, c0_n22_w46, c0_n22_w47, c0_n22_w48, c0_n22_w49, c0_n22_w50, c0_n22_w51, c0_n22_w52, c0_n22_w53, c0_n22_w54, c0_n22_w55, c0_n22_w56, c0_n22_w57, c0_n22_w58, c0_n22_w59, c0_n22_w60, c0_n22_w61, c0_n22_w62, c0_n22_w63, c0_n22_w64, c0_n22_w65, c0_n22_w66, c0_n22_w67, c0_n22_w68, c0_n22_w69, c0_n22_w70, c0_n22_w71, c0_n22_w72, c0_n22_w73, c0_n22_w74, c0_n22_w75, c0_n23_w1, c0_n23_w2, c0_n23_w3, c0_n23_w4, c0_n23_w5, c0_n23_w6, c0_n23_w7, c0_n23_w8, c0_n23_w9, c0_n23_w10, c0_n23_w11, c0_n23_w12, c0_n23_w13, c0_n23_w14, c0_n23_w15, c0_n23_w16, c0_n23_w17, c0_n23_w18, c0_n23_w19, c0_n23_w20, c0_n23_w21, c0_n23_w22, c0_n23_w23, c0_n23_w24, c0_n23_w25, c0_n23_w26, c0_n23_w27, c0_n23_w28, c0_n23_w29, c0_n23_w30, c0_n23_w31, c0_n23_w32, c0_n23_w33, c0_n23_w34, c0_n23_w35, c0_n23_w36, c0_n23_w37, c0_n23_w38, c0_n23_w39, c0_n23_w40, c0_n23_w41, c0_n23_w42, c0_n23_w43, c0_n23_w44, c0_n23_w45, c0_n23_w46, c0_n23_w47, c0_n23_w48, c0_n23_w49, c0_n23_w50, c0_n23_w51, c0_n23_w52, c0_n23_w53, c0_n23_w54, c0_n23_w55, c0_n23_w56, c0_n23_w57, c0_n23_w58, c0_n23_w59, c0_n23_w60, c0_n23_w61, c0_n23_w62, c0_n23_w63, c0_n23_w64, c0_n23_w65, c0_n23_w66, c0_n23_w67, c0_n23_w68, c0_n23_w69, c0_n23_w70, c0_n23_w71, c0_n23_w72, c0_n23_w73, c0_n23_w74, c0_n23_w75, c0_n24_w1, c0_n24_w2, c0_n24_w3, c0_n24_w4, c0_n24_w5, c0_n24_w6, c0_n24_w7, c0_n24_w8, c0_n24_w9, c0_n24_w10, c0_n24_w11, c0_n24_w12, c0_n24_w13, c0_n24_w14, c0_n24_w15, c0_n24_w16, c0_n24_w17, c0_n24_w18, c0_n24_w19, c0_n24_w20, c0_n24_w21, c0_n24_w22, c0_n24_w23, c0_n24_w24, c0_n24_w25, c0_n24_w26, c0_n24_w27, c0_n24_w28, c0_n24_w29, c0_n24_w30, c0_n24_w31, c0_n24_w32, c0_n24_w33, c0_n24_w34, c0_n24_w35, c0_n24_w36, c0_n24_w37, c0_n24_w38, c0_n24_w39, c0_n24_w40, c0_n24_w41, c0_n24_w42, c0_n24_w43, c0_n24_w44, c0_n24_w45, c0_n24_w46, c0_n24_w47, c0_n24_w48, c0_n24_w49, c0_n24_w50, c0_n24_w51, c0_n24_w52, c0_n24_w53, c0_n24_w54, c0_n24_w55, c0_n24_w56, c0_n24_w57, c0_n24_w58, c0_n24_w59, c0_n24_w60, c0_n24_w61, c0_n24_w62, c0_n24_w63, c0_n24_w64, c0_n24_w65, c0_n24_w66, c0_n24_w67, c0_n24_w68, c0_n24_w69, c0_n24_w70, c0_n24_w71, c0_n24_w72, c0_n24_w73, c0_n24_w74, c0_n24_w75, c0_n25_w1, c0_n25_w2, c0_n25_w3, c0_n25_w4, c0_n25_w5, c0_n25_w6, c0_n25_w7, c0_n25_w8, c0_n25_w9, c0_n25_w10, c0_n25_w11, c0_n25_w12, c0_n25_w13, c0_n25_w14, c0_n25_w15, c0_n25_w16, c0_n25_w17, c0_n25_w18, c0_n25_w19, c0_n25_w20, c0_n25_w21, c0_n25_w22, c0_n25_w23, c0_n25_w24, c0_n25_w25, c0_n25_w26, c0_n25_w27, c0_n25_w28, c0_n25_w29, c0_n25_w30, c0_n25_w31, c0_n25_w32, c0_n25_w33, c0_n25_w34, c0_n25_w35, c0_n25_w36, c0_n25_w37, c0_n25_w38, c0_n25_w39, c0_n25_w40, c0_n25_w41, c0_n25_w42, c0_n25_w43, c0_n25_w44, c0_n25_w45, c0_n25_w46, c0_n25_w47, c0_n25_w48, c0_n25_w49, c0_n25_w50, c0_n25_w51, c0_n25_w52, c0_n25_w53, c0_n25_w54, c0_n25_w55, c0_n25_w56, c0_n25_w57, c0_n25_w58, c0_n25_w59, c0_n25_w60, c0_n25_w61, c0_n25_w62, c0_n25_w63, c0_n25_w64, c0_n25_w65, c0_n25_w66, c0_n25_w67, c0_n25_w68, c0_n25_w69, c0_n25_w70, c0_n25_w71, c0_n25_w72, c0_n25_w73, c0_n25_w74, c0_n25_w75, c0_n26_w1, c0_n26_w2, c0_n26_w3, c0_n26_w4, c0_n26_w5, c0_n26_w6, c0_n26_w7, c0_n26_w8, c0_n26_w9, c0_n26_w10, c0_n26_w11, c0_n26_w12, c0_n26_w13, c0_n26_w14, c0_n26_w15, c0_n26_w16, c0_n26_w17, c0_n26_w18, c0_n26_w19, c0_n26_w20, c0_n26_w21, c0_n26_w22, c0_n26_w23, c0_n26_w24, c0_n26_w25, c0_n26_w26, c0_n26_w27, c0_n26_w28, c0_n26_w29, c0_n26_w30, c0_n26_w31, c0_n26_w32, c0_n26_w33, c0_n26_w34, c0_n26_w35, c0_n26_w36, c0_n26_w37, c0_n26_w38, c0_n26_w39, c0_n26_w40, c0_n26_w41, c0_n26_w42, c0_n26_w43, c0_n26_w44, c0_n26_w45, c0_n26_w46, c0_n26_w47, c0_n26_w48, c0_n26_w49, c0_n26_w50, c0_n26_w51, c0_n26_w52, c0_n26_w53, c0_n26_w54, c0_n26_w55, c0_n26_w56, c0_n26_w57, c0_n26_w58, c0_n26_w59, c0_n26_w60, c0_n26_w61, c0_n26_w62, c0_n26_w63, c0_n26_w64, c0_n26_w65, c0_n26_w66, c0_n26_w67, c0_n26_w68, c0_n26_w69, c0_n26_w70, c0_n26_w71, c0_n26_w72, c0_n26_w73, c0_n26_w74, c0_n26_w75, c0_n27_w1, c0_n27_w2, c0_n27_w3, c0_n27_w4, c0_n27_w5, c0_n27_w6, c0_n27_w7, c0_n27_w8, c0_n27_w9, c0_n27_w10, c0_n27_w11, c0_n27_w12, c0_n27_w13, c0_n27_w14, c0_n27_w15, c0_n27_w16, c0_n27_w17, c0_n27_w18, c0_n27_w19, c0_n27_w20, c0_n27_w21, c0_n27_w22, c0_n27_w23, c0_n27_w24, c0_n27_w25, c0_n27_w26, c0_n27_w27, c0_n27_w28, c0_n27_w29, c0_n27_w30, c0_n27_w31, c0_n27_w32, c0_n27_w33, c0_n27_w34, c0_n27_w35, c0_n27_w36, c0_n27_w37, c0_n27_w38, c0_n27_w39, c0_n27_w40, c0_n27_w41, c0_n27_w42, c0_n27_w43, c0_n27_w44, c0_n27_w45, c0_n27_w46, c0_n27_w47, c0_n27_w48, c0_n27_w49, c0_n27_w50, c0_n27_w51, c0_n27_w52, c0_n27_w53, c0_n27_w54, c0_n27_w55, c0_n27_w56, c0_n27_w57, c0_n27_w58, c0_n27_w59, c0_n27_w60, c0_n27_w61, c0_n27_w62, c0_n27_w63, c0_n27_w64, c0_n27_w65, c0_n27_w66, c0_n27_w67, c0_n27_w68, c0_n27_w69, c0_n27_w70, c0_n27_w71, c0_n27_w72, c0_n27_w73, c0_n27_w74, c0_n27_w75, c0_n28_w1, c0_n28_w2, c0_n28_w3, c0_n28_w4, c0_n28_w5, c0_n28_w6, c0_n28_w7, c0_n28_w8, c0_n28_w9, c0_n28_w10, c0_n28_w11, c0_n28_w12, c0_n28_w13, c0_n28_w14, c0_n28_w15, c0_n28_w16, c0_n28_w17, c0_n28_w18, c0_n28_w19, c0_n28_w20, c0_n28_w21, c0_n28_w22, c0_n28_w23, c0_n28_w24, c0_n28_w25, c0_n28_w26, c0_n28_w27, c0_n28_w28, c0_n28_w29, c0_n28_w30, c0_n28_w31, c0_n28_w32, c0_n28_w33, c0_n28_w34, c0_n28_w35, c0_n28_w36, c0_n28_w37, c0_n28_w38, c0_n28_w39, c0_n28_w40, c0_n28_w41, c0_n28_w42, c0_n28_w43, c0_n28_w44, c0_n28_w45, c0_n28_w46, c0_n28_w47, c0_n28_w48, c0_n28_w49, c0_n28_w50, c0_n28_w51, c0_n28_w52, c0_n28_w53, c0_n28_w54, c0_n28_w55, c0_n28_w56, c0_n28_w57, c0_n28_w58, c0_n28_w59, c0_n28_w60, c0_n28_w61, c0_n28_w62, c0_n28_w63, c0_n28_w64, c0_n28_w65, c0_n28_w66, c0_n28_w67, c0_n28_w68, c0_n28_w69, c0_n28_w70, c0_n28_w71, c0_n28_w72, c0_n28_w73, c0_n28_w74, c0_n28_w75, c0_n29_w1, c0_n29_w2, c0_n29_w3, c0_n29_w4, c0_n29_w5, c0_n29_w6, c0_n29_w7, c0_n29_w8, c0_n29_w9, c0_n29_w10, c0_n29_w11, c0_n29_w12, c0_n29_w13, c0_n29_w14, c0_n29_w15, c0_n29_w16, c0_n29_w17, c0_n29_w18, c0_n29_w19, c0_n29_w20, c0_n29_w21, c0_n29_w22, c0_n29_w23, c0_n29_w24, c0_n29_w25, c0_n29_w26, c0_n29_w27, c0_n29_w28, c0_n29_w29, c0_n29_w30, c0_n29_w31, c0_n29_w32, c0_n29_w33, c0_n29_w34, c0_n29_w35, c0_n29_w36, c0_n29_w37, c0_n29_w38, c0_n29_w39, c0_n29_w40, c0_n29_w41, c0_n29_w42, c0_n29_w43, c0_n29_w44, c0_n29_w45, c0_n29_w46, c0_n29_w47, c0_n29_w48, c0_n29_w49, c0_n29_w50, c0_n29_w51, c0_n29_w52, c0_n29_w53, c0_n29_w54, c0_n29_w55, c0_n29_w56, c0_n29_w57, c0_n29_w58, c0_n29_w59, c0_n29_w60, c0_n29_w61, c0_n29_w62, c0_n29_w63, c0_n29_w64, c0_n29_w65, c0_n29_w66, c0_n29_w67, c0_n29_w68, c0_n29_w69, c0_n29_w70, c0_n29_w71, c0_n29_w72, c0_n29_w73, c0_n29_w74, c0_n29_w75, c0_n30_w1, c0_n30_w2, c0_n30_w3, c0_n30_w4, c0_n30_w5, c0_n30_w6, c0_n30_w7, c0_n30_w8, c0_n30_w9, c0_n30_w10, c0_n30_w11, c0_n30_w12, c0_n30_w13, c0_n30_w14, c0_n30_w15, c0_n30_w16, c0_n30_w17, c0_n30_w18, c0_n30_w19, c0_n30_w20, c0_n30_w21, c0_n30_w22, c0_n30_w23, c0_n30_w24, c0_n30_w25, c0_n30_w26, c0_n30_w27, c0_n30_w28, c0_n30_w29, c0_n30_w30, c0_n30_w31, c0_n30_w32, c0_n30_w33, c0_n30_w34, c0_n30_w35, c0_n30_w36, c0_n30_w37, c0_n30_w38, c0_n30_w39, c0_n30_w40, c0_n30_w41, c0_n30_w42, c0_n30_w43, c0_n30_w44, c0_n30_w45, c0_n30_w46, c0_n30_w47, c0_n30_w48, c0_n30_w49, c0_n30_w50, c0_n30_w51, c0_n30_w52, c0_n30_w53, c0_n30_w54, c0_n30_w55, c0_n30_w56, c0_n30_w57, c0_n30_w58, c0_n30_w59, c0_n30_w60, c0_n30_w61, c0_n30_w62, c0_n30_w63, c0_n30_w64, c0_n30_w65, c0_n30_w66, c0_n30_w67, c0_n30_w68, c0_n30_w69, c0_n30_w70, c0_n30_w71, c0_n30_w72, c0_n30_w73, c0_n30_w74, c0_n30_w75, c0_n31_w1, c0_n31_w2, c0_n31_w3, c0_n31_w4, c0_n31_w5, c0_n31_w6, c0_n31_w7, c0_n31_w8, c0_n31_w9, c0_n31_w10, c0_n31_w11, c0_n31_w12, c0_n31_w13, c0_n31_w14, c0_n31_w15, c0_n31_w16, c0_n31_w17, c0_n31_w18, c0_n31_w19, c0_n31_w20, c0_n31_w21, c0_n31_w22, c0_n31_w23, c0_n31_w24, c0_n31_w25, c0_n31_w26, c0_n31_w27, c0_n31_w28, c0_n31_w29, c0_n31_w30, c0_n31_w31, c0_n31_w32, c0_n31_w33, c0_n31_w34, c0_n31_w35, c0_n31_w36, c0_n31_w37, c0_n31_w38, c0_n31_w39, c0_n31_w40, c0_n31_w41, c0_n31_w42, c0_n31_w43, c0_n31_w44, c0_n31_w45, c0_n31_w46, c0_n31_w47, c0_n31_w48, c0_n31_w49, c0_n31_w50, c0_n31_w51, c0_n31_w52, c0_n31_w53, c0_n31_w54, c0_n31_w55, c0_n31_w56, c0_n31_w57, c0_n31_w58, c0_n31_w59, c0_n31_w60, c0_n31_w61, c0_n31_w62, c0_n31_w63, c0_n31_w64, c0_n31_w65, c0_n31_w66, c0_n31_w67, c0_n31_w68, c0_n31_w69, c0_n31_w70, c0_n31_w71, c0_n31_w72, c0_n31_w73, c0_n31_w74, c0_n31_w75, c0_n32_w1, c0_n32_w2, c0_n32_w3, c0_n32_w4, c0_n32_w5, c0_n32_w6, c0_n32_w7, c0_n32_w8, c0_n32_w9, c0_n32_w10, c0_n32_w11, c0_n32_w12, c0_n32_w13, c0_n32_w14, c0_n32_w15, c0_n32_w16, c0_n32_w17, c0_n32_w18, c0_n32_w19, c0_n32_w20, c0_n32_w21, c0_n32_w22, c0_n32_w23, c0_n32_w24, c0_n32_w25, c0_n32_w26, c0_n32_w27, c0_n32_w28, c0_n32_w29, c0_n32_w30, c0_n32_w31, c0_n32_w32, c0_n32_w33, c0_n32_w34, c0_n32_w35, c0_n32_w36, c0_n32_w37, c0_n32_w38, c0_n32_w39, c0_n32_w40, c0_n32_w41, c0_n32_w42, c0_n32_w43, c0_n32_w44, c0_n32_w45, c0_n32_w46, c0_n32_w47, c0_n32_w48, c0_n32_w49, c0_n32_w50, c0_n32_w51, c0_n32_w52, c0_n32_w53, c0_n32_w54, c0_n32_w55, c0_n32_w56, c0_n32_w57, c0_n32_w58, c0_n32_w59, c0_n32_w60, c0_n32_w61, c0_n32_w62, c0_n32_w63, c0_n32_w64, c0_n32_w65, c0_n32_w66, c0_n32_w67, c0_n32_w68, c0_n32_w69, c0_n32_w70, c0_n32_w71, c0_n32_w72, c0_n32_w73, c0_n32_w74, c0_n32_w75, c0_n33_w1, c0_n33_w2, c0_n33_w3, c0_n33_w4, c0_n33_w5, c0_n33_w6, c0_n33_w7, c0_n33_w8, c0_n33_w9, c0_n33_w10, c0_n33_w11, c0_n33_w12, c0_n33_w13, c0_n33_w14, c0_n33_w15, c0_n33_w16, c0_n33_w17, c0_n33_w18, c0_n33_w19, c0_n33_w20, c0_n33_w21, c0_n33_w22, c0_n33_w23, c0_n33_w24, c0_n33_w25, c0_n33_w26, c0_n33_w27, c0_n33_w28, c0_n33_w29, c0_n33_w30, c0_n33_w31, c0_n33_w32, c0_n33_w33, c0_n33_w34, c0_n33_w35, c0_n33_w36, c0_n33_w37, c0_n33_w38, c0_n33_w39, c0_n33_w40, c0_n33_w41, c0_n33_w42, c0_n33_w43, c0_n33_w44, c0_n33_w45, c0_n33_w46, c0_n33_w47, c0_n33_w48, c0_n33_w49, c0_n33_w50, c0_n33_w51, c0_n33_w52, c0_n33_w53, c0_n33_w54, c0_n33_w55, c0_n33_w56, c0_n33_w57, c0_n33_w58, c0_n33_w59, c0_n33_w60, c0_n33_w61, c0_n33_w62, c0_n33_w63, c0_n33_w64, c0_n33_w65, c0_n33_w66, c0_n33_w67, c0_n33_w68, c0_n33_w69, c0_n33_w70, c0_n33_w71, c0_n33_w72, c0_n33_w73, c0_n33_w74, c0_n33_w75, c0_n34_w1, c0_n34_w2, c0_n34_w3, c0_n34_w4, c0_n34_w5, c0_n34_w6, c0_n34_w7, c0_n34_w8, c0_n34_w9, c0_n34_w10, c0_n34_w11, c0_n34_w12, c0_n34_w13, c0_n34_w14, c0_n34_w15, c0_n34_w16, c0_n34_w17, c0_n34_w18, c0_n34_w19, c0_n34_w20, c0_n34_w21, c0_n34_w22, c0_n34_w23, c0_n34_w24, c0_n34_w25, c0_n34_w26, c0_n34_w27, c0_n34_w28, c0_n34_w29, c0_n34_w30, c0_n34_w31, c0_n34_w32, c0_n34_w33, c0_n34_w34, c0_n34_w35, c0_n34_w36, c0_n34_w37, c0_n34_w38, c0_n34_w39, c0_n34_w40, c0_n34_w41, c0_n34_w42, c0_n34_w43, c0_n34_w44, c0_n34_w45, c0_n34_w46, c0_n34_w47, c0_n34_w48, c0_n34_w49, c0_n34_w50, c0_n34_w51, c0_n34_w52, c0_n34_w53, c0_n34_w54, c0_n34_w55, c0_n34_w56, c0_n34_w57, c0_n34_w58, c0_n34_w59, c0_n34_w60, c0_n34_w61, c0_n34_w62, c0_n34_w63, c0_n34_w64, c0_n34_w65, c0_n34_w66, c0_n34_w67, c0_n34_w68, c0_n34_w69, c0_n34_w70, c0_n34_w71, c0_n34_w72, c0_n34_w73, c0_n34_w74, c0_n34_w75, c0_n35_w1, c0_n35_w2, c0_n35_w3, c0_n35_w4, c0_n35_w5, c0_n35_w6, c0_n35_w7, c0_n35_w8, c0_n35_w9, c0_n35_w10, c0_n35_w11, c0_n35_w12, c0_n35_w13, c0_n35_w14, c0_n35_w15, c0_n35_w16, c0_n35_w17, c0_n35_w18, c0_n35_w19, c0_n35_w20, c0_n35_w21, c0_n35_w22, c0_n35_w23, c0_n35_w24, c0_n35_w25, c0_n35_w26, c0_n35_w27, c0_n35_w28, c0_n35_w29, c0_n35_w30, c0_n35_w31, c0_n35_w32, c0_n35_w33, c0_n35_w34, c0_n35_w35, c0_n35_w36, c0_n35_w37, c0_n35_w38, c0_n35_w39, c0_n35_w40, c0_n35_w41, c0_n35_w42, c0_n35_w43, c0_n35_w44, c0_n35_w45, c0_n35_w46, c0_n35_w47, c0_n35_w48, c0_n35_w49, c0_n35_w50, c0_n35_w51, c0_n35_w52, c0_n35_w53, c0_n35_w54, c0_n35_w55, c0_n35_w56, c0_n35_w57, c0_n35_w58, c0_n35_w59, c0_n35_w60, c0_n35_w61, c0_n35_w62, c0_n35_w63, c0_n35_w64, c0_n35_w65, c0_n35_w66, c0_n35_w67, c0_n35_w68, c0_n35_w69, c0_n35_w70, c0_n35_w71, c0_n35_w72, c0_n35_w73, c0_n35_w74, c0_n35_w75, c0_n36_w1, c0_n36_w2, c0_n36_w3, c0_n36_w4, c0_n36_w5, c0_n36_w6, c0_n36_w7, c0_n36_w8, c0_n36_w9, c0_n36_w10, c0_n36_w11, c0_n36_w12, c0_n36_w13, c0_n36_w14, c0_n36_w15, c0_n36_w16, c0_n36_w17, c0_n36_w18, c0_n36_w19, c0_n36_w20, c0_n36_w21, c0_n36_w22, c0_n36_w23, c0_n36_w24, c0_n36_w25, c0_n36_w26, c0_n36_w27, c0_n36_w28, c0_n36_w29, c0_n36_w30, c0_n36_w31, c0_n36_w32, c0_n36_w33, c0_n36_w34, c0_n36_w35, c0_n36_w36, c0_n36_w37, c0_n36_w38, c0_n36_w39, c0_n36_w40, c0_n36_w41, c0_n36_w42, c0_n36_w43, c0_n36_w44, c0_n36_w45, c0_n36_w46, c0_n36_w47, c0_n36_w48, c0_n36_w49, c0_n36_w50, c0_n36_w51, c0_n36_w52, c0_n36_w53, c0_n36_w54, c0_n36_w55, c0_n36_w56, c0_n36_w57, c0_n36_w58, c0_n36_w59, c0_n36_w60, c0_n36_w61, c0_n36_w62, c0_n36_w63, c0_n36_w64, c0_n36_w65, c0_n36_w66, c0_n36_w67, c0_n36_w68, c0_n36_w69, c0_n36_w70, c0_n36_w71, c0_n36_w72, c0_n36_w73, c0_n36_w74, c0_n36_w75, c0_n37_w1, c0_n37_w2, c0_n37_w3, c0_n37_w4, c0_n37_w5, c0_n37_w6, c0_n37_w7, c0_n37_w8, c0_n37_w9, c0_n37_w10, c0_n37_w11, c0_n37_w12, c0_n37_w13, c0_n37_w14, c0_n37_w15, c0_n37_w16, c0_n37_w17, c0_n37_w18, c0_n37_w19, c0_n37_w20, c0_n37_w21, c0_n37_w22, c0_n37_w23, c0_n37_w24, c0_n37_w25, c0_n37_w26, c0_n37_w27, c0_n37_w28, c0_n37_w29, c0_n37_w30, c0_n37_w31, c0_n37_w32, c0_n37_w33, c0_n37_w34, c0_n37_w35, c0_n37_w36, c0_n37_w37, c0_n37_w38, c0_n37_w39, c0_n37_w40, c0_n37_w41, c0_n37_w42, c0_n37_w43, c0_n37_w44, c0_n37_w45, c0_n37_w46, c0_n37_w47, c0_n37_w48, c0_n37_w49, c0_n37_w50, c0_n37_w51, c0_n37_w52, c0_n37_w53, c0_n37_w54, c0_n37_w55, c0_n37_w56, c0_n37_w57, c0_n37_w58, c0_n37_w59, c0_n37_w60, c0_n37_w61, c0_n37_w62, c0_n37_w63, c0_n37_w64, c0_n37_w65, c0_n37_w66, c0_n37_w67, c0_n37_w68, c0_n37_w69, c0_n37_w70, c0_n37_w71, c0_n37_w72, c0_n37_w73, c0_n37_w74, c0_n37_w75, c0_n38_w1, c0_n38_w2, c0_n38_w3, c0_n38_w4, c0_n38_w5, c0_n38_w6, c0_n38_w7, c0_n38_w8, c0_n38_w9, c0_n38_w10, c0_n38_w11, c0_n38_w12, c0_n38_w13, c0_n38_w14, c0_n38_w15, c0_n38_w16, c0_n38_w17, c0_n38_w18, c0_n38_w19, c0_n38_w20, c0_n38_w21, c0_n38_w22, c0_n38_w23, c0_n38_w24, c0_n38_w25, c0_n38_w26, c0_n38_w27, c0_n38_w28, c0_n38_w29, c0_n38_w30, c0_n38_w31, c0_n38_w32, c0_n38_w33, c0_n38_w34, c0_n38_w35, c0_n38_w36, c0_n38_w37, c0_n38_w38, c0_n38_w39, c0_n38_w40, c0_n38_w41, c0_n38_w42, c0_n38_w43, c0_n38_w44, c0_n38_w45, c0_n38_w46, c0_n38_w47, c0_n38_w48, c0_n38_w49, c0_n38_w50, c0_n38_w51, c0_n38_w52, c0_n38_w53, c0_n38_w54, c0_n38_w55, c0_n38_w56, c0_n38_w57, c0_n38_w58, c0_n38_w59, c0_n38_w60, c0_n38_w61, c0_n38_w62, c0_n38_w63, c0_n38_w64, c0_n38_w65, c0_n38_w66, c0_n38_w67, c0_n38_w68, c0_n38_w69, c0_n38_w70, c0_n38_w71, c0_n38_w72, c0_n38_w73, c0_n38_w74, c0_n38_w75, c0_n39_w1, c0_n39_w2, c0_n39_w3, c0_n39_w4, c0_n39_w5, c0_n39_w6, c0_n39_w7, c0_n39_w8, c0_n39_w9, c0_n39_w10, c0_n39_w11, c0_n39_w12, c0_n39_w13, c0_n39_w14, c0_n39_w15, c0_n39_w16, c0_n39_w17, c0_n39_w18, c0_n39_w19, c0_n39_w20, c0_n39_w21, c0_n39_w22, c0_n39_w23, c0_n39_w24, c0_n39_w25, c0_n39_w26, c0_n39_w27, c0_n39_w28, c0_n39_w29, c0_n39_w30, c0_n39_w31, c0_n39_w32, c0_n39_w33, c0_n39_w34, c0_n39_w35, c0_n39_w36, c0_n39_w37, c0_n39_w38, c0_n39_w39, c0_n39_w40, c0_n39_w41, c0_n39_w42, c0_n39_w43, c0_n39_w44, c0_n39_w45, c0_n39_w46, c0_n39_w47, c0_n39_w48, c0_n39_w49, c0_n39_w50, c0_n39_w51, c0_n39_w52, c0_n39_w53, c0_n39_w54, c0_n39_w55, c0_n39_w56, c0_n39_w57, c0_n39_w58, c0_n39_w59, c0_n39_w60, c0_n39_w61, c0_n39_w62, c0_n39_w63, c0_n39_w64, c0_n39_w65, c0_n39_w66, c0_n39_w67, c0_n39_w68, c0_n39_w69, c0_n39_w70, c0_n39_w71, c0_n39_w72, c0_n39_w73, c0_n39_w74, c0_n39_w75, c0_n40_w1, c0_n40_w2, c0_n40_w3, c0_n40_w4, c0_n40_w5, c0_n40_w6, c0_n40_w7, c0_n40_w8, c0_n40_w9, c0_n40_w10, c0_n40_w11, c0_n40_w12, c0_n40_w13, c0_n40_w14, c0_n40_w15, c0_n40_w16, c0_n40_w17, c0_n40_w18, c0_n40_w19, c0_n40_w20, c0_n40_w21, c0_n40_w22, c0_n40_w23, c0_n40_w24, c0_n40_w25, c0_n40_w26, c0_n40_w27, c0_n40_w28, c0_n40_w29, c0_n40_w30, c0_n40_w31, c0_n40_w32, c0_n40_w33, c0_n40_w34, c0_n40_w35, c0_n40_w36, c0_n40_w37, c0_n40_w38, c0_n40_w39, c0_n40_w40, c0_n40_w41, c0_n40_w42, c0_n40_w43, c0_n40_w44, c0_n40_w45, c0_n40_w46, c0_n40_w47, c0_n40_w48, c0_n40_w49, c0_n40_w50, c0_n40_w51, c0_n40_w52, c0_n40_w53, c0_n40_w54, c0_n40_w55, c0_n40_w56, c0_n40_w57, c0_n40_w58, c0_n40_w59, c0_n40_w60, c0_n40_w61, c0_n40_w62, c0_n40_w63, c0_n40_w64, c0_n40_w65, c0_n40_w66, c0_n40_w67, c0_n40_w68, c0_n40_w69, c0_n40_w70, c0_n40_w71, c0_n40_w72, c0_n40_w73, c0_n40_w74, c0_n40_w75, c0_n41_w1, c0_n41_w2, c0_n41_w3, c0_n41_w4, c0_n41_w5, c0_n41_w6, c0_n41_w7, c0_n41_w8, c0_n41_w9, c0_n41_w10, c0_n41_w11, c0_n41_w12, c0_n41_w13, c0_n41_w14, c0_n41_w15, c0_n41_w16, c0_n41_w17, c0_n41_w18, c0_n41_w19, c0_n41_w20, c0_n41_w21, c0_n41_w22, c0_n41_w23, c0_n41_w24, c0_n41_w25, c0_n41_w26, c0_n41_w27, c0_n41_w28, c0_n41_w29, c0_n41_w30, c0_n41_w31, c0_n41_w32, c0_n41_w33, c0_n41_w34, c0_n41_w35, c0_n41_w36, c0_n41_w37, c0_n41_w38, c0_n41_w39, c0_n41_w40, c0_n41_w41, c0_n41_w42, c0_n41_w43, c0_n41_w44, c0_n41_w45, c0_n41_w46, c0_n41_w47, c0_n41_w48, c0_n41_w49, c0_n41_w50, c0_n41_w51, c0_n41_w52, c0_n41_w53, c0_n41_w54, c0_n41_w55, c0_n41_w56, c0_n41_w57, c0_n41_w58, c0_n41_w59, c0_n41_w60, c0_n41_w61, c0_n41_w62, c0_n41_w63, c0_n41_w64, c0_n41_w65, c0_n41_w66, c0_n41_w67, c0_n41_w68, c0_n41_w69, c0_n41_w70, c0_n41_w71, c0_n41_w72, c0_n41_w73, c0_n41_w74, c0_n41_w75, c0_n42_w1, c0_n42_w2, c0_n42_w3, c0_n42_w4, c0_n42_w5, c0_n42_w6, c0_n42_w7, c0_n42_w8, c0_n42_w9, c0_n42_w10, c0_n42_w11, c0_n42_w12, c0_n42_w13, c0_n42_w14, c0_n42_w15, c0_n42_w16, c0_n42_w17, c0_n42_w18, c0_n42_w19, c0_n42_w20, c0_n42_w21, c0_n42_w22, c0_n42_w23, c0_n42_w24, c0_n42_w25, c0_n42_w26, c0_n42_w27, c0_n42_w28, c0_n42_w29, c0_n42_w30, c0_n42_w31, c0_n42_w32, c0_n42_w33, c0_n42_w34, c0_n42_w35, c0_n42_w36, c0_n42_w37, c0_n42_w38, c0_n42_w39, c0_n42_w40, c0_n42_w41, c0_n42_w42, c0_n42_w43, c0_n42_w44, c0_n42_w45, c0_n42_w46, c0_n42_w47, c0_n42_w48, c0_n42_w49, c0_n42_w50, c0_n42_w51, c0_n42_w52, c0_n42_w53, c0_n42_w54, c0_n42_w55, c0_n42_w56, c0_n42_w57, c0_n42_w58, c0_n42_w59, c0_n42_w60, c0_n42_w61, c0_n42_w62, c0_n42_w63, c0_n42_w64, c0_n42_w65, c0_n42_w66, c0_n42_w67, c0_n42_w68, c0_n42_w69, c0_n42_w70, c0_n42_w71, c0_n42_w72, c0_n42_w73, c0_n42_w74, c0_n42_w75, c0_n43_w1, c0_n43_w2, c0_n43_w3, c0_n43_w4, c0_n43_w5, c0_n43_w6, c0_n43_w7, c0_n43_w8, c0_n43_w9, c0_n43_w10, c0_n43_w11, c0_n43_w12, c0_n43_w13, c0_n43_w14, c0_n43_w15, c0_n43_w16, c0_n43_w17, c0_n43_w18, c0_n43_w19, c0_n43_w20, c0_n43_w21, c0_n43_w22, c0_n43_w23, c0_n43_w24, c0_n43_w25, c0_n43_w26, c0_n43_w27, c0_n43_w28, c0_n43_w29, c0_n43_w30, c0_n43_w31, c0_n43_w32, c0_n43_w33, c0_n43_w34, c0_n43_w35, c0_n43_w36, c0_n43_w37, c0_n43_w38, c0_n43_w39, c0_n43_w40, c0_n43_w41, c0_n43_w42, c0_n43_w43, c0_n43_w44, c0_n43_w45, c0_n43_w46, c0_n43_w47, c0_n43_w48, c0_n43_w49, c0_n43_w50, c0_n43_w51, c0_n43_w52, c0_n43_w53, c0_n43_w54, c0_n43_w55, c0_n43_w56, c0_n43_w57, c0_n43_w58, c0_n43_w59, c0_n43_w60, c0_n43_w61, c0_n43_w62, c0_n43_w63, c0_n43_w64, c0_n43_w65, c0_n43_w66, c0_n43_w67, c0_n43_w68, c0_n43_w69, c0_n43_w70, c0_n43_w71, c0_n43_w72, c0_n43_w73, c0_n43_w74, c0_n43_w75, c0_n44_w1, c0_n44_w2, c0_n44_w3, c0_n44_w4, c0_n44_w5, c0_n44_w6, c0_n44_w7, c0_n44_w8, c0_n44_w9, c0_n44_w10, c0_n44_w11, c0_n44_w12, c0_n44_w13, c0_n44_w14, c0_n44_w15, c0_n44_w16, c0_n44_w17, c0_n44_w18, c0_n44_w19, c0_n44_w20, c0_n44_w21, c0_n44_w22, c0_n44_w23, c0_n44_w24, c0_n44_w25, c0_n44_w26, c0_n44_w27, c0_n44_w28, c0_n44_w29, c0_n44_w30, c0_n44_w31, c0_n44_w32, c0_n44_w33, c0_n44_w34, c0_n44_w35, c0_n44_w36, c0_n44_w37, c0_n44_w38, c0_n44_w39, c0_n44_w40, c0_n44_w41, c0_n44_w42, c0_n44_w43, c0_n44_w44, c0_n44_w45, c0_n44_w46, c0_n44_w47, c0_n44_w48, c0_n44_w49, c0_n44_w50, c0_n44_w51, c0_n44_w52, c0_n44_w53, c0_n44_w54, c0_n44_w55, c0_n44_w56, c0_n44_w57, c0_n44_w58, c0_n44_w59, c0_n44_w60, c0_n44_w61, c0_n44_w62, c0_n44_w63, c0_n44_w64, c0_n44_w65, c0_n44_w66, c0_n44_w67, c0_n44_w68, c0_n44_w69, c0_n44_w70, c0_n44_w71, c0_n44_w72, c0_n44_w73, c0_n44_w74, c0_n44_w75, c0_n45_w1, c0_n45_w2, c0_n45_w3, c0_n45_w4, c0_n45_w5, c0_n45_w6, c0_n45_w7, c0_n45_w8, c0_n45_w9, c0_n45_w10, c0_n45_w11, c0_n45_w12, c0_n45_w13, c0_n45_w14, c0_n45_w15, c0_n45_w16, c0_n45_w17, c0_n45_w18, c0_n45_w19, c0_n45_w20, c0_n45_w21, c0_n45_w22, c0_n45_w23, c0_n45_w24, c0_n45_w25, c0_n45_w26, c0_n45_w27, c0_n45_w28, c0_n45_w29, c0_n45_w30, c0_n45_w31, c0_n45_w32, c0_n45_w33, c0_n45_w34, c0_n45_w35, c0_n45_w36, c0_n45_w37, c0_n45_w38, c0_n45_w39, c0_n45_w40, c0_n45_w41, c0_n45_w42, c0_n45_w43, c0_n45_w44, c0_n45_w45, c0_n45_w46, c0_n45_w47, c0_n45_w48, c0_n45_w49, c0_n45_w50, c0_n45_w51, c0_n45_w52, c0_n45_w53, c0_n45_w54, c0_n45_w55, c0_n45_w56, c0_n45_w57, c0_n45_w58, c0_n45_w59, c0_n45_w60, c0_n45_w61, c0_n45_w62, c0_n45_w63, c0_n45_w64, c0_n45_w65, c0_n45_w66, c0_n45_w67, c0_n45_w68, c0_n45_w69, c0_n45_w70, c0_n45_w71, c0_n45_w72, c0_n45_w73, c0_n45_w74, c0_n45_w75, c0_n46_w1, c0_n46_w2, c0_n46_w3, c0_n46_w4, c0_n46_w5, c0_n46_w6, c0_n46_w7, c0_n46_w8, c0_n46_w9, c0_n46_w10, c0_n46_w11, c0_n46_w12, c0_n46_w13, c0_n46_w14, c0_n46_w15, c0_n46_w16, c0_n46_w17, c0_n46_w18, c0_n46_w19, c0_n46_w20, c0_n46_w21, c0_n46_w22, c0_n46_w23, c0_n46_w24, c0_n46_w25, c0_n46_w26, c0_n46_w27, c0_n46_w28, c0_n46_w29, c0_n46_w30, c0_n46_w31, c0_n46_w32, c0_n46_w33, c0_n46_w34, c0_n46_w35, c0_n46_w36, c0_n46_w37, c0_n46_w38, c0_n46_w39, c0_n46_w40, c0_n46_w41, c0_n46_w42, c0_n46_w43, c0_n46_w44, c0_n46_w45, c0_n46_w46, c0_n46_w47, c0_n46_w48, c0_n46_w49, c0_n46_w50, c0_n46_w51, c0_n46_w52, c0_n46_w53, c0_n46_w54, c0_n46_w55, c0_n46_w56, c0_n46_w57, c0_n46_w58, c0_n46_w59, c0_n46_w60, c0_n46_w61, c0_n46_w62, c0_n46_w63, c0_n46_w64, c0_n46_w65, c0_n46_w66, c0_n46_w67, c0_n46_w68, c0_n46_w69, c0_n46_w70, c0_n46_w71, c0_n46_w72, c0_n46_w73, c0_n46_w74, c0_n46_w75, c0_n47_w1, c0_n47_w2, c0_n47_w3, c0_n47_w4, c0_n47_w5, c0_n47_w6, c0_n47_w7, c0_n47_w8, c0_n47_w9, c0_n47_w10, c0_n47_w11, c0_n47_w12, c0_n47_w13, c0_n47_w14, c0_n47_w15, c0_n47_w16, c0_n47_w17, c0_n47_w18, c0_n47_w19, c0_n47_w20, c0_n47_w21, c0_n47_w22, c0_n47_w23, c0_n47_w24, c0_n47_w25, c0_n47_w26, c0_n47_w27, c0_n47_w28, c0_n47_w29, c0_n47_w30, c0_n47_w31, c0_n47_w32, c0_n47_w33, c0_n47_w34, c0_n47_w35, c0_n47_w36, c0_n47_w37, c0_n47_w38, c0_n47_w39, c0_n47_w40, c0_n47_w41, c0_n47_w42, c0_n47_w43, c0_n47_w44, c0_n47_w45, c0_n47_w46, c0_n47_w47, c0_n47_w48, c0_n47_w49, c0_n47_w50, c0_n47_w51, c0_n47_w52, c0_n47_w53, c0_n47_w54, c0_n47_w55, c0_n47_w56, c0_n47_w57, c0_n47_w58, c0_n47_w59, c0_n47_w60, c0_n47_w61, c0_n47_w62, c0_n47_w63, c0_n47_w64, c0_n47_w65, c0_n47_w66, c0_n47_w67, c0_n47_w68, c0_n47_w69, c0_n47_w70, c0_n47_w71, c0_n47_w72, c0_n47_w73, c0_n47_w74, c0_n47_w75, c0_n48_w1, c0_n48_w2, c0_n48_w3, c0_n48_w4, c0_n48_w5, c0_n48_w6, c0_n48_w7, c0_n48_w8, c0_n48_w9, c0_n48_w10, c0_n48_w11, c0_n48_w12, c0_n48_w13, c0_n48_w14, c0_n48_w15, c0_n48_w16, c0_n48_w17, c0_n48_w18, c0_n48_w19, c0_n48_w20, c0_n48_w21, c0_n48_w22, c0_n48_w23, c0_n48_w24, c0_n48_w25, c0_n48_w26, c0_n48_w27, c0_n48_w28, c0_n48_w29, c0_n48_w30, c0_n48_w31, c0_n48_w32, c0_n48_w33, c0_n48_w34, c0_n48_w35, c0_n48_w36, c0_n48_w37, c0_n48_w38, c0_n48_w39, c0_n48_w40, c0_n48_w41, c0_n48_w42, c0_n48_w43, c0_n48_w44, c0_n48_w45, c0_n48_w46, c0_n48_w47, c0_n48_w48, c0_n48_w49, c0_n48_w50, c0_n48_w51, c0_n48_w52, c0_n48_w53, c0_n48_w54, c0_n48_w55, c0_n48_w56, c0_n48_w57, c0_n48_w58, c0_n48_w59, c0_n48_w60, c0_n48_w61, c0_n48_w62, c0_n48_w63, c0_n48_w64, c0_n48_w65, c0_n48_w66, c0_n48_w67, c0_n48_w68, c0_n48_w69, c0_n48_w70, c0_n48_w71, c0_n48_w72, c0_n48_w73, c0_n48_w74, c0_n48_w75, c0_n49_w1, c0_n49_w2, c0_n49_w3, c0_n49_w4, c0_n49_w5, c0_n49_w6, c0_n49_w7, c0_n49_w8, c0_n49_w9, c0_n49_w10, c0_n49_w11, c0_n49_w12, c0_n49_w13, c0_n49_w14, c0_n49_w15, c0_n49_w16, c0_n49_w17, c0_n49_w18, c0_n49_w19, c0_n49_w20, c0_n49_w21, c0_n49_w22, c0_n49_w23, c0_n49_w24, c0_n49_w25, c0_n49_w26, c0_n49_w27, c0_n49_w28, c0_n49_w29, c0_n49_w30, c0_n49_w31, c0_n49_w32, c0_n49_w33, c0_n49_w34, c0_n49_w35, c0_n49_w36, c0_n49_w37, c0_n49_w38, c0_n49_w39, c0_n49_w40, c0_n49_w41, c0_n49_w42, c0_n49_w43, c0_n49_w44, c0_n49_w45, c0_n49_w46, c0_n49_w47, c0_n49_w48, c0_n49_w49, c0_n49_w50, c0_n49_w51, c0_n49_w52, c0_n49_w53, c0_n49_w54, c0_n49_w55, c0_n49_w56, c0_n49_w57, c0_n49_w58, c0_n49_w59, c0_n49_w60, c0_n49_w61, c0_n49_w62, c0_n49_w63, c0_n49_w64, c0_n49_w65, c0_n49_w66, c0_n49_w67, c0_n49_w68, c0_n49_w69, c0_n49_w70, c0_n49_w71, c0_n49_w72, c0_n49_w73, c0_n49_w74, c0_n49_w75, c0_n50_w1, c0_n50_w2, c0_n50_w3, c0_n50_w4, c0_n50_w5, c0_n50_w6, c0_n50_w7, c0_n50_w8, c0_n50_w9, c0_n50_w10, c0_n50_w11, c0_n50_w12, c0_n50_w13, c0_n50_w14, c0_n50_w15, c0_n50_w16, c0_n50_w17, c0_n50_w18, c0_n50_w19, c0_n50_w20, c0_n50_w21, c0_n50_w22, c0_n50_w23, c0_n50_w24, c0_n50_w25, c0_n50_w26, c0_n50_w27, c0_n50_w28, c0_n50_w29, c0_n50_w30, c0_n50_w31, c0_n50_w32, c0_n50_w33, c0_n50_w34, c0_n50_w35, c0_n50_w36, c0_n50_w37, c0_n50_w38, c0_n50_w39, c0_n50_w40, c0_n50_w41, c0_n50_w42, c0_n50_w43, c0_n50_w44, c0_n50_w45, c0_n50_w46, c0_n50_w47, c0_n50_w48, c0_n50_w49, c0_n50_w50, c0_n50_w51, c0_n50_w52, c0_n50_w53, c0_n50_w54, c0_n50_w55, c0_n50_w56, c0_n50_w57, c0_n50_w58, c0_n50_w59, c0_n50_w60, c0_n50_w61, c0_n50_w62, c0_n50_w63, c0_n50_w64, c0_n50_w65, c0_n50_w66, c0_n50_w67, c0_n50_w68, c0_n50_w69, c0_n50_w70, c0_n50_w71, c0_n50_w72, c0_n50_w73, c0_n50_w74, c0_n50_w75, c0_n51_w1, c0_n51_w2, c0_n51_w3, c0_n51_w4, c0_n51_w5, c0_n51_w6, c0_n51_w7, c0_n51_w8, c0_n51_w9, c0_n51_w10, c0_n51_w11, c0_n51_w12, c0_n51_w13, c0_n51_w14, c0_n51_w15, c0_n51_w16, c0_n51_w17, c0_n51_w18, c0_n51_w19, c0_n51_w20, c0_n51_w21, c0_n51_w22, c0_n51_w23, c0_n51_w24, c0_n51_w25, c0_n51_w26, c0_n51_w27, c0_n51_w28, c0_n51_w29, c0_n51_w30, c0_n51_w31, c0_n51_w32, c0_n51_w33, c0_n51_w34, c0_n51_w35, c0_n51_w36, c0_n51_w37, c0_n51_w38, c0_n51_w39, c0_n51_w40, c0_n51_w41, c0_n51_w42, c0_n51_w43, c0_n51_w44, c0_n51_w45, c0_n51_w46, c0_n51_w47, c0_n51_w48, c0_n51_w49, c0_n51_w50, c0_n51_w51, c0_n51_w52, c0_n51_w53, c0_n51_w54, c0_n51_w55, c0_n51_w56, c0_n51_w57, c0_n51_w58, c0_n51_w59, c0_n51_w60, c0_n51_w61, c0_n51_w62, c0_n51_w63, c0_n51_w64, c0_n51_w65, c0_n51_w66, c0_n51_w67, c0_n51_w68, c0_n51_w69, c0_n51_w70, c0_n51_w71, c0_n51_w72, c0_n51_w73, c0_n51_w74, c0_n51_w75, c0_n52_w1, c0_n52_w2, c0_n52_w3, c0_n52_w4, c0_n52_w5, c0_n52_w6, c0_n52_w7, c0_n52_w8, c0_n52_w9, c0_n52_w10, c0_n52_w11, c0_n52_w12, c0_n52_w13, c0_n52_w14, c0_n52_w15, c0_n52_w16, c0_n52_w17, c0_n52_w18, c0_n52_w19, c0_n52_w20, c0_n52_w21, c0_n52_w22, c0_n52_w23, c0_n52_w24, c0_n52_w25, c0_n52_w26, c0_n52_w27, c0_n52_w28, c0_n52_w29, c0_n52_w30, c0_n52_w31, c0_n52_w32, c0_n52_w33, c0_n52_w34, c0_n52_w35, c0_n52_w36, c0_n52_w37, c0_n52_w38, c0_n52_w39, c0_n52_w40, c0_n52_w41, c0_n52_w42, c0_n52_w43, c0_n52_w44, c0_n52_w45, c0_n52_w46, c0_n52_w47, c0_n52_w48, c0_n52_w49, c0_n52_w50, c0_n52_w51, c0_n52_w52, c0_n52_w53, c0_n52_w54, c0_n52_w55, c0_n52_w56, c0_n52_w57, c0_n52_w58, c0_n52_w59, c0_n52_w60, c0_n52_w61, c0_n52_w62, c0_n52_w63, c0_n52_w64, c0_n52_w65, c0_n52_w66, c0_n52_w67, c0_n52_w68, c0_n52_w69, c0_n52_w70, c0_n52_w71, c0_n52_w72, c0_n52_w73, c0_n52_w74, c0_n52_w75, c0_n53_w1, c0_n53_w2, c0_n53_w3, c0_n53_w4, c0_n53_w5, c0_n53_w6, c0_n53_w7, c0_n53_w8, c0_n53_w9, c0_n53_w10, c0_n53_w11, c0_n53_w12, c0_n53_w13, c0_n53_w14, c0_n53_w15, c0_n53_w16, c0_n53_w17, c0_n53_w18, c0_n53_w19, c0_n53_w20, c0_n53_w21, c0_n53_w22, c0_n53_w23, c0_n53_w24, c0_n53_w25, c0_n53_w26, c0_n53_w27, c0_n53_w28, c0_n53_w29, c0_n53_w30, c0_n53_w31, c0_n53_w32, c0_n53_w33, c0_n53_w34, c0_n53_w35, c0_n53_w36, c0_n53_w37, c0_n53_w38, c0_n53_w39, c0_n53_w40, c0_n53_w41, c0_n53_w42, c0_n53_w43, c0_n53_w44, c0_n53_w45, c0_n53_w46, c0_n53_w47, c0_n53_w48, c0_n53_w49, c0_n53_w50, c0_n53_w51, c0_n53_w52, c0_n53_w53, c0_n53_w54, c0_n53_w55, c0_n53_w56, c0_n53_w57, c0_n53_w58, c0_n53_w59, c0_n53_w60, c0_n53_w61, c0_n53_w62, c0_n53_w63, c0_n53_w64, c0_n53_w65, c0_n53_w66, c0_n53_w67, c0_n53_w68, c0_n53_w69, c0_n53_w70, c0_n53_w71, c0_n53_w72, c0_n53_w73, c0_n53_w74, c0_n53_w75, c0_n54_w1, c0_n54_w2, c0_n54_w3, c0_n54_w4, c0_n54_w5, c0_n54_w6, c0_n54_w7, c0_n54_w8, c0_n54_w9, c0_n54_w10, c0_n54_w11, c0_n54_w12, c0_n54_w13, c0_n54_w14, c0_n54_w15, c0_n54_w16, c0_n54_w17, c0_n54_w18, c0_n54_w19, c0_n54_w20, c0_n54_w21, c0_n54_w22, c0_n54_w23, c0_n54_w24, c0_n54_w25, c0_n54_w26, c0_n54_w27, c0_n54_w28, c0_n54_w29, c0_n54_w30, c0_n54_w31, c0_n54_w32, c0_n54_w33, c0_n54_w34, c0_n54_w35, c0_n54_w36, c0_n54_w37, c0_n54_w38, c0_n54_w39, c0_n54_w40, c0_n54_w41, c0_n54_w42, c0_n54_w43, c0_n54_w44, c0_n54_w45, c0_n54_w46, c0_n54_w47, c0_n54_w48, c0_n54_w49, c0_n54_w50, c0_n54_w51, c0_n54_w52, c0_n54_w53, c0_n54_w54, c0_n54_w55, c0_n54_w56, c0_n54_w57, c0_n54_w58, c0_n54_w59, c0_n54_w60, c0_n54_w61, c0_n54_w62, c0_n54_w63, c0_n54_w64, c0_n54_w65, c0_n54_w66, c0_n54_w67, c0_n54_w68, c0_n54_w69, c0_n54_w70, c0_n54_w71, c0_n54_w72, c0_n54_w73, c0_n54_w74, c0_n54_w75, c0_n55_w1, c0_n55_w2, c0_n55_w3, c0_n55_w4, c0_n55_w5, c0_n55_w6, c0_n55_w7, c0_n55_w8, c0_n55_w9, c0_n55_w10, c0_n55_w11, c0_n55_w12, c0_n55_w13, c0_n55_w14, c0_n55_w15, c0_n55_w16, c0_n55_w17, c0_n55_w18, c0_n55_w19, c0_n55_w20, c0_n55_w21, c0_n55_w22, c0_n55_w23, c0_n55_w24, c0_n55_w25, c0_n55_w26, c0_n55_w27, c0_n55_w28, c0_n55_w29, c0_n55_w30, c0_n55_w31, c0_n55_w32, c0_n55_w33, c0_n55_w34, c0_n55_w35, c0_n55_w36, c0_n55_w37, c0_n55_w38, c0_n55_w39, c0_n55_w40, c0_n55_w41, c0_n55_w42, c0_n55_w43, c0_n55_w44, c0_n55_w45, c0_n55_w46, c0_n55_w47, c0_n55_w48, c0_n55_w49, c0_n55_w50, c0_n55_w51, c0_n55_w52, c0_n55_w53, c0_n55_w54, c0_n55_w55, c0_n55_w56, c0_n55_w57, c0_n55_w58, c0_n55_w59, c0_n55_w60, c0_n55_w61, c0_n55_w62, c0_n55_w63, c0_n55_w64, c0_n55_w65, c0_n55_w66, c0_n55_w67, c0_n55_w68, c0_n55_w69, c0_n55_w70, c0_n55_w71, c0_n55_w72, c0_n55_w73, c0_n55_w74, c0_n55_w75, c0_n56_w1, c0_n56_w2, c0_n56_w3, c0_n56_w4, c0_n56_w5, c0_n56_w6, c0_n56_w7, c0_n56_w8, c0_n56_w9, c0_n56_w10, c0_n56_w11, c0_n56_w12, c0_n56_w13, c0_n56_w14, c0_n56_w15, c0_n56_w16, c0_n56_w17, c0_n56_w18, c0_n56_w19, c0_n56_w20, c0_n56_w21, c0_n56_w22, c0_n56_w23, c0_n56_w24, c0_n56_w25, c0_n56_w26, c0_n56_w27, c0_n56_w28, c0_n56_w29, c0_n56_w30, c0_n56_w31, c0_n56_w32, c0_n56_w33, c0_n56_w34, c0_n56_w35, c0_n56_w36, c0_n56_w37, c0_n56_w38, c0_n56_w39, c0_n56_w40, c0_n56_w41, c0_n56_w42, c0_n56_w43, c0_n56_w44, c0_n56_w45, c0_n56_w46, c0_n56_w47, c0_n56_w48, c0_n56_w49, c0_n56_w50, c0_n56_w51, c0_n56_w52, c0_n56_w53, c0_n56_w54, c0_n56_w55, c0_n56_w56, c0_n56_w57, c0_n56_w58, c0_n56_w59, c0_n56_w60, c0_n56_w61, c0_n56_w62, c0_n56_w63, c0_n56_w64, c0_n56_w65, c0_n56_w66, c0_n56_w67, c0_n56_w68, c0_n56_w69, c0_n56_w70, c0_n56_w71, c0_n56_w72, c0_n56_w73, c0_n56_w74, c0_n56_w75, c0_n57_w1, c0_n57_w2, c0_n57_w3, c0_n57_w4, c0_n57_w5, c0_n57_w6, c0_n57_w7, c0_n57_w8, c0_n57_w9, c0_n57_w10, c0_n57_w11, c0_n57_w12, c0_n57_w13, c0_n57_w14, c0_n57_w15, c0_n57_w16, c0_n57_w17, c0_n57_w18, c0_n57_w19, c0_n57_w20, c0_n57_w21, c0_n57_w22, c0_n57_w23, c0_n57_w24, c0_n57_w25, c0_n57_w26, c0_n57_w27, c0_n57_w28, c0_n57_w29, c0_n57_w30, c0_n57_w31, c0_n57_w32, c0_n57_w33, c0_n57_w34, c0_n57_w35, c0_n57_w36, c0_n57_w37, c0_n57_w38, c0_n57_w39, c0_n57_w40, c0_n57_w41, c0_n57_w42, c0_n57_w43, c0_n57_w44, c0_n57_w45, c0_n57_w46, c0_n57_w47, c0_n57_w48, c0_n57_w49, c0_n57_w50, c0_n57_w51, c0_n57_w52, c0_n57_w53, c0_n57_w54, c0_n57_w55, c0_n57_w56, c0_n57_w57, c0_n57_w58, c0_n57_w59, c0_n57_w60, c0_n57_w61, c0_n57_w62, c0_n57_w63, c0_n57_w64, c0_n57_w65, c0_n57_w66, c0_n57_w67, c0_n57_w68, c0_n57_w69, c0_n57_w70, c0_n57_w71, c0_n57_w72, c0_n57_w73, c0_n57_w74, c0_n57_w75, c0_n58_w1, c0_n58_w2, c0_n58_w3, c0_n58_w4, c0_n58_w5, c0_n58_w6, c0_n58_w7, c0_n58_w8, c0_n58_w9, c0_n58_w10, c0_n58_w11, c0_n58_w12, c0_n58_w13, c0_n58_w14, c0_n58_w15, c0_n58_w16, c0_n58_w17, c0_n58_w18, c0_n58_w19, c0_n58_w20, c0_n58_w21, c0_n58_w22, c0_n58_w23, c0_n58_w24, c0_n58_w25, c0_n58_w26, c0_n58_w27, c0_n58_w28, c0_n58_w29, c0_n58_w30, c0_n58_w31, c0_n58_w32, c0_n58_w33, c0_n58_w34, c0_n58_w35, c0_n58_w36, c0_n58_w37, c0_n58_w38, c0_n58_w39, c0_n58_w40, c0_n58_w41, c0_n58_w42, c0_n58_w43, c0_n58_w44, c0_n58_w45, c0_n58_w46, c0_n58_w47, c0_n58_w48, c0_n58_w49, c0_n58_w50, c0_n58_w51, c0_n58_w52, c0_n58_w53, c0_n58_w54, c0_n58_w55, c0_n58_w56, c0_n58_w57, c0_n58_w58, c0_n58_w59, c0_n58_w60, c0_n58_w61, c0_n58_w62, c0_n58_w63, c0_n58_w64, c0_n58_w65, c0_n58_w66, c0_n58_w67, c0_n58_w68, c0_n58_w69, c0_n58_w70, c0_n58_w71, c0_n58_w72, c0_n58_w73, c0_n58_w74, c0_n58_w75, c0_n59_w1, c0_n59_w2, c0_n59_w3, c0_n59_w4, c0_n59_w5, c0_n59_w6, c0_n59_w7, c0_n59_w8, c0_n59_w9, c0_n59_w10, c0_n59_w11, c0_n59_w12, c0_n59_w13, c0_n59_w14, c0_n59_w15, c0_n59_w16, c0_n59_w17, c0_n59_w18, c0_n59_w19, c0_n59_w20, c0_n59_w21, c0_n59_w22, c0_n59_w23, c0_n59_w24, c0_n59_w25, c0_n59_w26, c0_n59_w27, c0_n59_w28, c0_n59_w29, c0_n59_w30, c0_n59_w31, c0_n59_w32, c0_n59_w33, c0_n59_w34, c0_n59_w35, c0_n59_w36, c0_n59_w37, c0_n59_w38, c0_n59_w39, c0_n59_w40, c0_n59_w41, c0_n59_w42, c0_n59_w43, c0_n59_w44, c0_n59_w45, c0_n59_w46, c0_n59_w47, c0_n59_w48, c0_n59_w49, c0_n59_w50, c0_n59_w51, c0_n59_w52, c0_n59_w53, c0_n59_w54, c0_n59_w55, c0_n59_w56, c0_n59_w57, c0_n59_w58, c0_n59_w59, c0_n59_w60, c0_n59_w61, c0_n59_w62, c0_n59_w63, c0_n59_w64, c0_n59_w65, c0_n59_w66, c0_n59_w67, c0_n59_w68, c0_n59_w69, c0_n59_w70, c0_n59_w71, c0_n59_w72, c0_n59_w73, c0_n59_w74, c0_n59_w75, c0_n60_w1, c0_n60_w2, c0_n60_w3, c0_n60_w4, c0_n60_w5, c0_n60_w6, c0_n60_w7, c0_n60_w8, c0_n60_w9, c0_n60_w10, c0_n60_w11, c0_n60_w12, c0_n60_w13, c0_n60_w14, c0_n60_w15, c0_n60_w16, c0_n60_w17, c0_n60_w18, c0_n60_w19, c0_n60_w20, c0_n60_w21, c0_n60_w22, c0_n60_w23, c0_n60_w24, c0_n60_w25, c0_n60_w26, c0_n60_w27, c0_n60_w28, c0_n60_w29, c0_n60_w30, c0_n60_w31, c0_n60_w32, c0_n60_w33, c0_n60_w34, c0_n60_w35, c0_n60_w36, c0_n60_w37, c0_n60_w38, c0_n60_w39, c0_n60_w40, c0_n60_w41, c0_n60_w42, c0_n60_w43, c0_n60_w44, c0_n60_w45, c0_n60_w46, c0_n60_w47, c0_n60_w48, c0_n60_w49, c0_n60_w50, c0_n60_w51, c0_n60_w52, c0_n60_w53, c0_n60_w54, c0_n60_w55, c0_n60_w56, c0_n60_w57, c0_n60_w58, c0_n60_w59, c0_n60_w60, c0_n60_w61, c0_n60_w62, c0_n60_w63, c0_n60_w64, c0_n60_w65, c0_n60_w66, c0_n60_w67, c0_n60_w68, c0_n60_w69, c0_n60_w70, c0_n60_w71, c0_n60_w72, c0_n60_w73, c0_n60_w74, c0_n60_w75, c0_n61_w1, c0_n61_w2, c0_n61_w3, c0_n61_w4, c0_n61_w5, c0_n61_w6, c0_n61_w7, c0_n61_w8, c0_n61_w9, c0_n61_w10, c0_n61_w11, c0_n61_w12, c0_n61_w13, c0_n61_w14, c0_n61_w15, c0_n61_w16, c0_n61_w17, c0_n61_w18, c0_n61_w19, c0_n61_w20, c0_n61_w21, c0_n61_w22, c0_n61_w23, c0_n61_w24, c0_n61_w25, c0_n61_w26, c0_n61_w27, c0_n61_w28, c0_n61_w29, c0_n61_w30, c0_n61_w31, c0_n61_w32, c0_n61_w33, c0_n61_w34, c0_n61_w35, c0_n61_w36, c0_n61_w37, c0_n61_w38, c0_n61_w39, c0_n61_w40, c0_n61_w41, c0_n61_w42, c0_n61_w43, c0_n61_w44, c0_n61_w45, c0_n61_w46, c0_n61_w47, c0_n61_w48, c0_n61_w49, c0_n61_w50, c0_n61_w51, c0_n61_w52, c0_n61_w53, c0_n61_w54, c0_n61_w55, c0_n61_w56, c0_n61_w57, c0_n61_w58, c0_n61_w59, c0_n61_w60, c0_n61_w61, c0_n61_w62, c0_n61_w63, c0_n61_w64, c0_n61_w65, c0_n61_w66, c0_n61_w67, c0_n61_w68, c0_n61_w69, c0_n61_w70, c0_n61_w71, c0_n61_w72, c0_n61_w73, c0_n61_w74, c0_n61_w75, c0_n62_w1, c0_n62_w2, c0_n62_w3, c0_n62_w4, c0_n62_w5, c0_n62_w6, c0_n62_w7, c0_n62_w8, c0_n62_w9, c0_n62_w10, c0_n62_w11, c0_n62_w12, c0_n62_w13, c0_n62_w14, c0_n62_w15, c0_n62_w16, c0_n62_w17, c0_n62_w18, c0_n62_w19, c0_n62_w20, c0_n62_w21, c0_n62_w22, c0_n62_w23, c0_n62_w24, c0_n62_w25, c0_n62_w26, c0_n62_w27, c0_n62_w28, c0_n62_w29, c0_n62_w30, c0_n62_w31, c0_n62_w32, c0_n62_w33, c0_n62_w34, c0_n62_w35, c0_n62_w36, c0_n62_w37, c0_n62_w38, c0_n62_w39, c0_n62_w40, c0_n62_w41, c0_n62_w42, c0_n62_w43, c0_n62_w44, c0_n62_w45, c0_n62_w46, c0_n62_w47, c0_n62_w48, c0_n62_w49, c0_n62_w50, c0_n62_w51, c0_n62_w52, c0_n62_w53, c0_n62_w54, c0_n62_w55, c0_n62_w56, c0_n62_w57, c0_n62_w58, c0_n62_w59, c0_n62_w60, c0_n62_w61, c0_n62_w62, c0_n62_w63, c0_n62_w64, c0_n62_w65, c0_n62_w66, c0_n62_w67, c0_n62_w68, c0_n62_w69, c0_n62_w70, c0_n62_w71, c0_n62_w72, c0_n62_w73, c0_n62_w74, c0_n62_w75, c0_n63_w1, c0_n63_w2, c0_n63_w3, c0_n63_w4, c0_n63_w5, c0_n63_w6, c0_n63_w7, c0_n63_w8, c0_n63_w9, c0_n63_w10, c0_n63_w11, c0_n63_w12, c0_n63_w13, c0_n63_w14, c0_n63_w15, c0_n63_w16, c0_n63_w17, c0_n63_w18, c0_n63_w19, c0_n63_w20, c0_n63_w21, c0_n63_w22, c0_n63_w23, c0_n63_w24, c0_n63_w25, c0_n63_w26, c0_n63_w27, c0_n63_w28, c0_n63_w29, c0_n63_w30, c0_n63_w31, c0_n63_w32, c0_n63_w33, c0_n63_w34, c0_n63_w35, c0_n63_w36, c0_n63_w37, c0_n63_w38, c0_n63_w39, c0_n63_w40, c0_n63_w41, c0_n63_w42, c0_n63_w43, c0_n63_w44, c0_n63_w45, c0_n63_w46, c0_n63_w47, c0_n63_w48, c0_n63_w49, c0_n63_w50, c0_n63_w51, c0_n63_w52, c0_n63_w53, c0_n63_w54, c0_n63_w55, c0_n63_w56, c0_n63_w57, c0_n63_w58, c0_n63_w59, c0_n63_w60, c0_n63_w61, c0_n63_w62, c0_n63_w63, c0_n63_w64, c0_n63_w65, c0_n63_w66, c0_n63_w67, c0_n63_w68, c0_n63_w69, c0_n63_w70, c0_n63_w71, c0_n63_w72, c0_n63_w73, c0_n63_w74, c0_n63_w75, c0_n64_w1, c0_n64_w2, c0_n64_w3, c0_n64_w4, c0_n64_w5, c0_n64_w6, c0_n64_w7, c0_n64_w8, c0_n64_w9, c0_n64_w10, c0_n64_w11, c0_n64_w12, c0_n64_w13, c0_n64_w14, c0_n64_w15, c0_n64_w16, c0_n64_w17, c0_n64_w18, c0_n64_w19, c0_n64_w20, c0_n64_w21, c0_n64_w22, c0_n64_w23, c0_n64_w24, c0_n64_w25, c0_n64_w26, c0_n64_w27, c0_n64_w28, c0_n64_w29, c0_n64_w30, c0_n64_w31, c0_n64_w32, c0_n64_w33, c0_n64_w34, c0_n64_w35, c0_n64_w36, c0_n64_w37, c0_n64_w38, c0_n64_w39, c0_n64_w40, c0_n64_w41, c0_n64_w42, c0_n64_w43, c0_n64_w44, c0_n64_w45, c0_n64_w46, c0_n64_w47, c0_n64_w48, c0_n64_w49, c0_n64_w50, c0_n64_w51, c0_n64_w52, c0_n64_w53, c0_n64_w54, c0_n64_w55, c0_n64_w56, c0_n64_w57, c0_n64_w58, c0_n64_w59, c0_n64_w60, c0_n64_w61, c0_n64_w62, c0_n64_w63, c0_n64_w64, c0_n64_w65, c0_n64_w66, c0_n64_w67, c0_n64_w68, c0_n64_w69, c0_n64_w70, c0_n64_w71, c0_n64_w72, c0_n64_w73, c0_n64_w74, c0_n64_w75, c0_n65_w1, c0_n65_w2, c0_n65_w3, c0_n65_w4, c0_n65_w5, c0_n65_w6, c0_n65_w7, c0_n65_w8, c0_n65_w9, c0_n65_w10, c0_n65_w11, c0_n65_w12, c0_n65_w13, c0_n65_w14, c0_n65_w15, c0_n65_w16, c0_n65_w17, c0_n65_w18, c0_n65_w19, c0_n65_w20, c0_n65_w21, c0_n65_w22, c0_n65_w23, c0_n65_w24, c0_n65_w25, c0_n65_w26, c0_n65_w27, c0_n65_w28, c0_n65_w29, c0_n65_w30, c0_n65_w31, c0_n65_w32, c0_n65_w33, c0_n65_w34, c0_n65_w35, c0_n65_w36, c0_n65_w37, c0_n65_w38, c0_n65_w39, c0_n65_w40, c0_n65_w41, c0_n65_w42, c0_n65_w43, c0_n65_w44, c0_n65_w45, c0_n65_w46, c0_n65_w47, c0_n65_w48, c0_n65_w49, c0_n65_w50, c0_n65_w51, c0_n65_w52, c0_n65_w53, c0_n65_w54, c0_n65_w55, c0_n65_w56, c0_n65_w57, c0_n65_w58, c0_n65_w59, c0_n65_w60, c0_n65_w61, c0_n65_w62, c0_n65_w63, c0_n65_w64, c0_n65_w65, c0_n65_w66, c0_n65_w67, c0_n65_w68, c0_n65_w69, c0_n65_w70, c0_n65_w71, c0_n65_w72, c0_n65_w73, c0_n65_w74, c0_n65_w75, c0_n66_w1, c0_n66_w2, c0_n66_w3, c0_n66_w4, c0_n66_w5, c0_n66_w6, c0_n66_w7, c0_n66_w8, c0_n66_w9, c0_n66_w10, c0_n66_w11, c0_n66_w12, c0_n66_w13, c0_n66_w14, c0_n66_w15, c0_n66_w16, c0_n66_w17, c0_n66_w18, c0_n66_w19, c0_n66_w20, c0_n66_w21, c0_n66_w22, c0_n66_w23, c0_n66_w24, c0_n66_w25, c0_n66_w26, c0_n66_w27, c0_n66_w28, c0_n66_w29, c0_n66_w30, c0_n66_w31, c0_n66_w32, c0_n66_w33, c0_n66_w34, c0_n66_w35, c0_n66_w36, c0_n66_w37, c0_n66_w38, c0_n66_w39, c0_n66_w40, c0_n66_w41, c0_n66_w42, c0_n66_w43, c0_n66_w44, c0_n66_w45, c0_n66_w46, c0_n66_w47, c0_n66_w48, c0_n66_w49, c0_n66_w50, c0_n66_w51, c0_n66_w52, c0_n66_w53, c0_n66_w54, c0_n66_w55, c0_n66_w56, c0_n66_w57, c0_n66_w58, c0_n66_w59, c0_n66_w60, c0_n66_w61, c0_n66_w62, c0_n66_w63, c0_n66_w64, c0_n66_w65, c0_n66_w66, c0_n66_w67, c0_n66_w68, c0_n66_w69, c0_n66_w70, c0_n66_w71, c0_n66_w72, c0_n66_w73, c0_n66_w74, c0_n66_w75, c0_n67_w1, c0_n67_w2, c0_n67_w3, c0_n67_w4, c0_n67_w5, c0_n67_w6, c0_n67_w7, c0_n67_w8, c0_n67_w9, c0_n67_w10, c0_n67_w11, c0_n67_w12, c0_n67_w13, c0_n67_w14, c0_n67_w15, c0_n67_w16, c0_n67_w17, c0_n67_w18, c0_n67_w19, c0_n67_w20, c0_n67_w21, c0_n67_w22, c0_n67_w23, c0_n67_w24, c0_n67_w25, c0_n67_w26, c0_n67_w27, c0_n67_w28, c0_n67_w29, c0_n67_w30, c0_n67_w31, c0_n67_w32, c0_n67_w33, c0_n67_w34, c0_n67_w35, c0_n67_w36, c0_n67_w37, c0_n67_w38, c0_n67_w39, c0_n67_w40, c0_n67_w41, c0_n67_w42, c0_n67_w43, c0_n67_w44, c0_n67_w45, c0_n67_w46, c0_n67_w47, c0_n67_w48, c0_n67_w49, c0_n67_w50, c0_n67_w51, c0_n67_w52, c0_n67_w53, c0_n67_w54, c0_n67_w55, c0_n67_w56, c0_n67_w57, c0_n67_w58, c0_n67_w59, c0_n67_w60, c0_n67_w61, c0_n67_w62, c0_n67_w63, c0_n67_w64, c0_n67_w65, c0_n67_w66, c0_n67_w67, c0_n67_w68, c0_n67_w69, c0_n67_w70, c0_n67_w71, c0_n67_w72, c0_n67_w73, c0_n67_w74, c0_n67_w75, c0_n68_w1, c0_n68_w2, c0_n68_w3, c0_n68_w4, c0_n68_w5, c0_n68_w6, c0_n68_w7, c0_n68_w8, c0_n68_w9, c0_n68_w10, c0_n68_w11, c0_n68_w12, c0_n68_w13, c0_n68_w14, c0_n68_w15, c0_n68_w16, c0_n68_w17, c0_n68_w18, c0_n68_w19, c0_n68_w20, c0_n68_w21, c0_n68_w22, c0_n68_w23, c0_n68_w24, c0_n68_w25, c0_n68_w26, c0_n68_w27, c0_n68_w28, c0_n68_w29, c0_n68_w30, c0_n68_w31, c0_n68_w32, c0_n68_w33, c0_n68_w34, c0_n68_w35, c0_n68_w36, c0_n68_w37, c0_n68_w38, c0_n68_w39, c0_n68_w40, c0_n68_w41, c0_n68_w42, c0_n68_w43, c0_n68_w44, c0_n68_w45, c0_n68_w46, c0_n68_w47, c0_n68_w48, c0_n68_w49, c0_n68_w50, c0_n68_w51, c0_n68_w52, c0_n68_w53, c0_n68_w54, c0_n68_w55, c0_n68_w56, c0_n68_w57, c0_n68_w58, c0_n68_w59, c0_n68_w60, c0_n68_w61, c0_n68_w62, c0_n68_w63, c0_n68_w64, c0_n68_w65, c0_n68_w66, c0_n68_w67, c0_n68_w68, c0_n68_w69, c0_n68_w70, c0_n68_w71, c0_n68_w72, c0_n68_w73, c0_n68_w74, c0_n68_w75, c0_n69_w1, c0_n69_w2, c0_n69_w3, c0_n69_w4, c0_n69_w5, c0_n69_w6, c0_n69_w7, c0_n69_w8, c0_n69_w9, c0_n69_w10, c0_n69_w11, c0_n69_w12, c0_n69_w13, c0_n69_w14, c0_n69_w15, c0_n69_w16, c0_n69_w17, c0_n69_w18, c0_n69_w19, c0_n69_w20, c0_n69_w21, c0_n69_w22, c0_n69_w23, c0_n69_w24, c0_n69_w25, c0_n69_w26, c0_n69_w27, c0_n69_w28, c0_n69_w29, c0_n69_w30, c0_n69_w31, c0_n69_w32, c0_n69_w33, c0_n69_w34, c0_n69_w35, c0_n69_w36, c0_n69_w37, c0_n69_w38, c0_n69_w39, c0_n69_w40, c0_n69_w41, c0_n69_w42, c0_n69_w43, c0_n69_w44, c0_n69_w45, c0_n69_w46, c0_n69_w47, c0_n69_w48, c0_n69_w49, c0_n69_w50, c0_n69_w51, c0_n69_w52, c0_n69_w53, c0_n69_w54, c0_n69_w55, c0_n69_w56, c0_n69_w57, c0_n69_w58, c0_n69_w59, c0_n69_w60, c0_n69_w61, c0_n69_w62, c0_n69_w63, c0_n69_w64, c0_n69_w65, c0_n69_w66, c0_n69_w67, c0_n69_w68, c0_n69_w69, c0_n69_w70, c0_n69_w71, c0_n69_w72, c0_n69_w73, c0_n69_w74, c0_n69_w75, c0_n70_w1, c0_n70_w2, c0_n70_w3, c0_n70_w4, c0_n70_w5, c0_n70_w6, c0_n70_w7, c0_n70_w8, c0_n70_w9, c0_n70_w10, c0_n70_w11, c0_n70_w12, c0_n70_w13, c0_n70_w14, c0_n70_w15, c0_n70_w16, c0_n70_w17, c0_n70_w18, c0_n70_w19, c0_n70_w20, c0_n70_w21, c0_n70_w22, c0_n70_w23, c0_n70_w24, c0_n70_w25, c0_n70_w26, c0_n70_w27, c0_n70_w28, c0_n70_w29, c0_n70_w30, c0_n70_w31, c0_n70_w32, c0_n70_w33, c0_n70_w34, c0_n70_w35, c0_n70_w36, c0_n70_w37, c0_n70_w38, c0_n70_w39, c0_n70_w40, c0_n70_w41, c0_n70_w42, c0_n70_w43, c0_n70_w44, c0_n70_w45, c0_n70_w46, c0_n70_w47, c0_n70_w48, c0_n70_w49, c0_n70_w50, c0_n70_w51, c0_n70_w52, c0_n70_w53, c0_n70_w54, c0_n70_w55, c0_n70_w56, c0_n70_w57, c0_n70_w58, c0_n70_w59, c0_n70_w60, c0_n70_w61, c0_n70_w62, c0_n70_w63, c0_n70_w64, c0_n70_w65, c0_n70_w66, c0_n70_w67, c0_n70_w68, c0_n70_w69, c0_n70_w70, c0_n70_w71, c0_n70_w72, c0_n70_w73, c0_n70_w74, c0_n70_w75, c0_n71_w1, c0_n71_w2, c0_n71_w3, c0_n71_w4, c0_n71_w5, c0_n71_w6, c0_n71_w7, c0_n71_w8, c0_n71_w9, c0_n71_w10, c0_n71_w11, c0_n71_w12, c0_n71_w13, c0_n71_w14, c0_n71_w15, c0_n71_w16, c0_n71_w17, c0_n71_w18, c0_n71_w19, c0_n71_w20, c0_n71_w21, c0_n71_w22, c0_n71_w23, c0_n71_w24, c0_n71_w25, c0_n71_w26, c0_n71_w27, c0_n71_w28, c0_n71_w29, c0_n71_w30, c0_n71_w31, c0_n71_w32, c0_n71_w33, c0_n71_w34, c0_n71_w35, c0_n71_w36, c0_n71_w37, c0_n71_w38, c0_n71_w39, c0_n71_w40, c0_n71_w41, c0_n71_w42, c0_n71_w43, c0_n71_w44, c0_n71_w45, c0_n71_w46, c0_n71_w47, c0_n71_w48, c0_n71_w49, c0_n71_w50, c0_n71_w51, c0_n71_w52, c0_n71_w53, c0_n71_w54, c0_n71_w55, c0_n71_w56, c0_n71_w57, c0_n71_w58, c0_n71_w59, c0_n71_w60, c0_n71_w61, c0_n71_w62, c0_n71_w63, c0_n71_w64, c0_n71_w65, c0_n71_w66, c0_n71_w67, c0_n71_w68, c0_n71_w69, c0_n71_w70, c0_n71_w71, c0_n71_w72, c0_n71_w73, c0_n71_w74, c0_n71_w75, c0_n72_w1, c0_n72_w2, c0_n72_w3, c0_n72_w4, c0_n72_w5, c0_n72_w6, c0_n72_w7, c0_n72_w8, c0_n72_w9, c0_n72_w10, c0_n72_w11, c0_n72_w12, c0_n72_w13, c0_n72_w14, c0_n72_w15, c0_n72_w16, c0_n72_w17, c0_n72_w18, c0_n72_w19, c0_n72_w20, c0_n72_w21, c0_n72_w22, c0_n72_w23, c0_n72_w24, c0_n72_w25, c0_n72_w26, c0_n72_w27, c0_n72_w28, c0_n72_w29, c0_n72_w30, c0_n72_w31, c0_n72_w32, c0_n72_w33, c0_n72_w34, c0_n72_w35, c0_n72_w36, c0_n72_w37, c0_n72_w38, c0_n72_w39, c0_n72_w40, c0_n72_w41, c0_n72_w42, c0_n72_w43, c0_n72_w44, c0_n72_w45, c0_n72_w46, c0_n72_w47, c0_n72_w48, c0_n72_w49, c0_n72_w50, c0_n72_w51, c0_n72_w52, c0_n72_w53, c0_n72_w54, c0_n72_w55, c0_n72_w56, c0_n72_w57, c0_n72_w58, c0_n72_w59, c0_n72_w60, c0_n72_w61, c0_n72_w62, c0_n72_w63, c0_n72_w64, c0_n72_w65, c0_n72_w66, c0_n72_w67, c0_n72_w68, c0_n72_w69, c0_n72_w70, c0_n72_w71, c0_n72_w72, c0_n72_w73, c0_n72_w74, c0_n72_w75, c0_n73_w1, c0_n73_w2, c0_n73_w3, c0_n73_w4, c0_n73_w5, c0_n73_w6, c0_n73_w7, c0_n73_w8, c0_n73_w9, c0_n73_w10, c0_n73_w11, c0_n73_w12, c0_n73_w13, c0_n73_w14, c0_n73_w15, c0_n73_w16, c0_n73_w17, c0_n73_w18, c0_n73_w19, c0_n73_w20, c0_n73_w21, c0_n73_w22, c0_n73_w23, c0_n73_w24, c0_n73_w25, c0_n73_w26, c0_n73_w27, c0_n73_w28, c0_n73_w29, c0_n73_w30, c0_n73_w31, c0_n73_w32, c0_n73_w33, c0_n73_w34, c0_n73_w35, c0_n73_w36, c0_n73_w37, c0_n73_w38, c0_n73_w39, c0_n73_w40, c0_n73_w41, c0_n73_w42, c0_n73_w43, c0_n73_w44, c0_n73_w45, c0_n73_w46, c0_n73_w47, c0_n73_w48, c0_n73_w49, c0_n73_w50, c0_n73_w51, c0_n73_w52, c0_n73_w53, c0_n73_w54, c0_n73_w55, c0_n73_w56, c0_n73_w57, c0_n73_w58, c0_n73_w59, c0_n73_w60, c0_n73_w61, c0_n73_w62, c0_n73_w63, c0_n73_w64, c0_n73_w65, c0_n73_w66, c0_n73_w67, c0_n73_w68, c0_n73_w69, c0_n73_w70, c0_n73_w71, c0_n73_w72, c0_n73_w73, c0_n73_w74, c0_n73_w75, c0_n74_w1, c0_n74_w2, c0_n74_w3, c0_n74_w4, c0_n74_w5, c0_n74_w6, c0_n74_w7, c0_n74_w8, c0_n74_w9, c0_n74_w10, c0_n74_w11, c0_n74_w12, c0_n74_w13, c0_n74_w14, c0_n74_w15, c0_n74_w16, c0_n74_w17, c0_n74_w18, c0_n74_w19, c0_n74_w20, c0_n74_w21, c0_n74_w22, c0_n74_w23, c0_n74_w24, c0_n74_w25, c0_n74_w26, c0_n74_w27, c0_n74_w28, c0_n74_w29, c0_n74_w30, c0_n74_w31, c0_n74_w32, c0_n74_w33, c0_n74_w34, c0_n74_w35, c0_n74_w36, c0_n74_w37, c0_n74_w38, c0_n74_w39, c0_n74_w40, c0_n74_w41, c0_n74_w42, c0_n74_w43, c0_n74_w44, c0_n74_w45, c0_n74_w46, c0_n74_w47, c0_n74_w48, c0_n74_w49, c0_n74_w50, c0_n74_w51, c0_n74_w52, c0_n74_w53, c0_n74_w54, c0_n74_w55, c0_n74_w56, c0_n74_w57, c0_n74_w58, c0_n74_w59, c0_n74_w60, c0_n74_w61, c0_n74_w62, c0_n74_w63, c0_n74_w64, c0_n74_w65, c0_n74_w66, c0_n74_w67, c0_n74_w68, c0_n74_w69, c0_n74_w70, c0_n74_w71, c0_n74_w72, c0_n74_w73, c0_n74_w74, c0_n74_w75, c0_n75_w1, c0_n75_w2, c0_n75_w3, c0_n75_w4, c0_n75_w5, c0_n75_w6, c0_n75_w7, c0_n75_w8, c0_n75_w9, c0_n75_w10, c0_n75_w11, c0_n75_w12, c0_n75_w13, c0_n75_w14, c0_n75_w15, c0_n75_w16, c0_n75_w17, c0_n75_w18, c0_n75_w19, c0_n75_w20, c0_n75_w21, c0_n75_w22, c0_n75_w23, c0_n75_w24, c0_n75_w25, c0_n75_w26, c0_n75_w27, c0_n75_w28, c0_n75_w29, c0_n75_w30, c0_n75_w31, c0_n75_w32, c0_n75_w33, c0_n75_w34, c0_n75_w35, c0_n75_w36, c0_n75_w37, c0_n75_w38, c0_n75_w39, c0_n75_w40, c0_n75_w41, c0_n75_w42, c0_n75_w43, c0_n75_w44, c0_n75_w45, c0_n75_w46, c0_n75_w47, c0_n75_w48, c0_n75_w49, c0_n75_w50, c0_n75_w51, c0_n75_w52, c0_n75_w53, c0_n75_w54, c0_n75_w55, c0_n75_w56, c0_n75_w57, c0_n75_w58, c0_n75_w59, c0_n75_w60, c0_n75_w61, c0_n75_w62, c0_n75_w63, c0_n75_w64, c0_n75_w65, c0_n75_w66, c0_n75_w67, c0_n75_w68, c0_n75_w69, c0_n75_w70, c0_n75_w71, c0_n75_w72, c0_n75_w73, c0_n75_w74, c0_n75_w75, c0_n76_w1, c0_n76_w2, c0_n76_w3, c0_n76_w4, c0_n76_w5, c0_n76_w6, c0_n76_w7, c0_n76_w8, c0_n76_w9, c0_n76_w10, c0_n76_w11, c0_n76_w12, c0_n76_w13, c0_n76_w14, c0_n76_w15, c0_n76_w16, c0_n76_w17, c0_n76_w18, c0_n76_w19, c0_n76_w20, c0_n76_w21, c0_n76_w22, c0_n76_w23, c0_n76_w24, c0_n76_w25, c0_n76_w26, c0_n76_w27, c0_n76_w28, c0_n76_w29, c0_n76_w30, c0_n76_w31, c0_n76_w32, c0_n76_w33, c0_n76_w34, c0_n76_w35, c0_n76_w36, c0_n76_w37, c0_n76_w38, c0_n76_w39, c0_n76_w40, c0_n76_w41, c0_n76_w42, c0_n76_w43, c0_n76_w44, c0_n76_w45, c0_n76_w46, c0_n76_w47, c0_n76_w48, c0_n76_w49, c0_n76_w50, c0_n76_w51, c0_n76_w52, c0_n76_w53, c0_n76_w54, c0_n76_w55, c0_n76_w56, c0_n76_w57, c0_n76_w58, c0_n76_w59, c0_n76_w60, c0_n76_w61, c0_n76_w62, c0_n76_w63, c0_n76_w64, c0_n76_w65, c0_n76_w66, c0_n76_w67, c0_n76_w68, c0_n76_w69, c0_n76_w70, c0_n76_w71, c0_n76_w72, c0_n76_w73, c0_n76_w74, c0_n76_w75, c0_n77_w1, c0_n77_w2, c0_n77_w3, c0_n77_w4, c0_n77_w5, c0_n77_w6, c0_n77_w7, c0_n77_w8, c0_n77_w9, c0_n77_w10, c0_n77_w11, c0_n77_w12, c0_n77_w13, c0_n77_w14, c0_n77_w15, c0_n77_w16, c0_n77_w17, c0_n77_w18, c0_n77_w19, c0_n77_w20, c0_n77_w21, c0_n77_w22, c0_n77_w23, c0_n77_w24, c0_n77_w25, c0_n77_w26, c0_n77_w27, c0_n77_w28, c0_n77_w29, c0_n77_w30, c0_n77_w31, c0_n77_w32, c0_n77_w33, c0_n77_w34, c0_n77_w35, c0_n77_w36, c0_n77_w37, c0_n77_w38, c0_n77_w39, c0_n77_w40, c0_n77_w41, c0_n77_w42, c0_n77_w43, c0_n77_w44, c0_n77_w45, c0_n77_w46, c0_n77_w47, c0_n77_w48, c0_n77_w49, c0_n77_w50, c0_n77_w51, c0_n77_w52, c0_n77_w53, c0_n77_w54, c0_n77_w55, c0_n77_w56, c0_n77_w57, c0_n77_w58, c0_n77_w59, c0_n77_w60, c0_n77_w61, c0_n77_w62, c0_n77_w63, c0_n77_w64, c0_n77_w65, c0_n77_w66, c0_n77_w67, c0_n77_w68, c0_n77_w69, c0_n77_w70, c0_n77_w71, c0_n77_w72, c0_n77_w73, c0_n77_w74, c0_n77_w75, c0_n78_w1, c0_n78_w2, c0_n78_w3, c0_n78_w4, c0_n78_w5, c0_n78_w6, c0_n78_w7, c0_n78_w8, c0_n78_w9, c0_n78_w10, c0_n78_w11, c0_n78_w12, c0_n78_w13, c0_n78_w14, c0_n78_w15, c0_n78_w16, c0_n78_w17, c0_n78_w18, c0_n78_w19, c0_n78_w20, c0_n78_w21, c0_n78_w22, c0_n78_w23, c0_n78_w24, c0_n78_w25, c0_n78_w26, c0_n78_w27, c0_n78_w28, c0_n78_w29, c0_n78_w30, c0_n78_w31, c0_n78_w32, c0_n78_w33, c0_n78_w34, c0_n78_w35, c0_n78_w36, c0_n78_w37, c0_n78_w38, c0_n78_w39, c0_n78_w40, c0_n78_w41, c0_n78_w42, c0_n78_w43, c0_n78_w44, c0_n78_w45, c0_n78_w46, c0_n78_w47, c0_n78_w48, c0_n78_w49, c0_n78_w50, c0_n78_w51, c0_n78_w52, c0_n78_w53, c0_n78_w54, c0_n78_w55, c0_n78_w56, c0_n78_w57, c0_n78_w58, c0_n78_w59, c0_n78_w60, c0_n78_w61, c0_n78_w62, c0_n78_w63, c0_n78_w64, c0_n78_w65, c0_n78_w66, c0_n78_w67, c0_n78_w68, c0_n78_w69, c0_n78_w70, c0_n78_w71, c0_n78_w72, c0_n78_w73, c0_n78_w74, c0_n78_w75, c0_n79_w1, c0_n79_w2, c0_n79_w3, c0_n79_w4, c0_n79_w5, c0_n79_w6, c0_n79_w7, c0_n79_w8, c0_n79_w9, c0_n79_w10, c0_n79_w11, c0_n79_w12, c0_n79_w13, c0_n79_w14, c0_n79_w15, c0_n79_w16, c0_n79_w17, c0_n79_w18, c0_n79_w19, c0_n79_w20, c0_n79_w21, c0_n79_w22, c0_n79_w23, c0_n79_w24, c0_n79_w25, c0_n79_w26, c0_n79_w27, c0_n79_w28, c0_n79_w29, c0_n79_w30, c0_n79_w31, c0_n79_w32, c0_n79_w33, c0_n79_w34, c0_n79_w35, c0_n79_w36, c0_n79_w37, c0_n79_w38, c0_n79_w39, c0_n79_w40, c0_n79_w41, c0_n79_w42, c0_n79_w43, c0_n79_w44, c0_n79_w45, c0_n79_w46, c0_n79_w47, c0_n79_w48, c0_n79_w49, c0_n79_w50, c0_n79_w51, c0_n79_w52, c0_n79_w53, c0_n79_w54, c0_n79_w55, c0_n79_w56, c0_n79_w57, c0_n79_w58, c0_n79_w59, c0_n79_w60, c0_n79_w61, c0_n79_w62, c0_n79_w63, c0_n79_w64, c0_n79_w65, c0_n79_w66, c0_n79_w67, c0_n79_w68, c0_n79_w69, c0_n79_w70, c0_n79_w71, c0_n79_w72, c0_n79_w73, c0_n79_w74, c0_n79_w75, c0_n80_w1, c0_n80_w2, c0_n80_w3, c0_n80_w4, c0_n80_w5, c0_n80_w6, c0_n80_w7, c0_n80_w8, c0_n80_w9, c0_n80_w10, c0_n80_w11, c0_n80_w12, c0_n80_w13, c0_n80_w14, c0_n80_w15, c0_n80_w16, c0_n80_w17, c0_n80_w18, c0_n80_w19, c0_n80_w20, c0_n80_w21, c0_n80_w22, c0_n80_w23, c0_n80_w24, c0_n80_w25, c0_n80_w26, c0_n80_w27, c0_n80_w28, c0_n80_w29, c0_n80_w30, c0_n80_w31, c0_n80_w32, c0_n80_w33, c0_n80_w34, c0_n80_w35, c0_n80_w36, c0_n80_w37, c0_n80_w38, c0_n80_w39, c0_n80_w40, c0_n80_w41, c0_n80_w42, c0_n80_w43, c0_n80_w44, c0_n80_w45, c0_n80_w46, c0_n80_w47, c0_n80_w48, c0_n80_w49, c0_n80_w50, c0_n80_w51, c0_n80_w52, c0_n80_w53, c0_n80_w54, c0_n80_w55, c0_n80_w56, c0_n80_w57, c0_n80_w58, c0_n80_w59, c0_n80_w60, c0_n80_w61, c0_n80_w62, c0_n80_w63, c0_n80_w64, c0_n80_w65, c0_n80_w66, c0_n80_w67, c0_n80_w68, c0_n80_w69, c0_n80_w70, c0_n80_w71, c0_n80_w72, c0_n80_w73, c0_n80_w74, c0_n80_w75, c0_n81_w1, c0_n81_w2, c0_n81_w3, c0_n81_w4, c0_n81_w5, c0_n81_w6, c0_n81_w7, c0_n81_w8, c0_n81_w9, c0_n81_w10, c0_n81_w11, c0_n81_w12, c0_n81_w13, c0_n81_w14, c0_n81_w15, c0_n81_w16, c0_n81_w17, c0_n81_w18, c0_n81_w19, c0_n81_w20, c0_n81_w21, c0_n81_w22, c0_n81_w23, c0_n81_w24, c0_n81_w25, c0_n81_w26, c0_n81_w27, c0_n81_w28, c0_n81_w29, c0_n81_w30, c0_n81_w31, c0_n81_w32, c0_n81_w33, c0_n81_w34, c0_n81_w35, c0_n81_w36, c0_n81_w37, c0_n81_w38, c0_n81_w39, c0_n81_w40, c0_n81_w41, c0_n81_w42, c0_n81_w43, c0_n81_w44, c0_n81_w45, c0_n81_w46, c0_n81_w47, c0_n81_w48, c0_n81_w49, c0_n81_w50, c0_n81_w51, c0_n81_w52, c0_n81_w53, c0_n81_w54, c0_n81_w55, c0_n81_w56, c0_n81_w57, c0_n81_w58, c0_n81_w59, c0_n81_w60, c0_n81_w61, c0_n81_w62, c0_n81_w63, c0_n81_w64, c0_n81_w65, c0_n81_w66, c0_n81_w67, c0_n81_w68, c0_n81_w69, c0_n81_w70, c0_n81_w71, c0_n81_w72, c0_n81_w73, c0_n81_w74, c0_n81_w75, c0_n82_w1, c0_n82_w2, c0_n82_w3, c0_n82_w4, c0_n82_w5, c0_n82_w6, c0_n82_w7, c0_n82_w8, c0_n82_w9, c0_n82_w10, c0_n82_w11, c0_n82_w12, c0_n82_w13, c0_n82_w14, c0_n82_w15, c0_n82_w16, c0_n82_w17, c0_n82_w18, c0_n82_w19, c0_n82_w20, c0_n82_w21, c0_n82_w22, c0_n82_w23, c0_n82_w24, c0_n82_w25, c0_n82_w26, c0_n82_w27, c0_n82_w28, c0_n82_w29, c0_n82_w30, c0_n82_w31, c0_n82_w32, c0_n82_w33, c0_n82_w34, c0_n82_w35, c0_n82_w36, c0_n82_w37, c0_n82_w38, c0_n82_w39, c0_n82_w40, c0_n82_w41, c0_n82_w42, c0_n82_w43, c0_n82_w44, c0_n82_w45, c0_n82_w46, c0_n82_w47, c0_n82_w48, c0_n82_w49, c0_n82_w50, c0_n82_w51, c0_n82_w52, c0_n82_w53, c0_n82_w54, c0_n82_w55, c0_n82_w56, c0_n82_w57, c0_n82_w58, c0_n82_w59, c0_n82_w60, c0_n82_w61, c0_n82_w62, c0_n82_w63, c0_n82_w64, c0_n82_w65, c0_n82_w66, c0_n82_w67, c0_n82_w68, c0_n82_w69, c0_n82_w70, c0_n82_w71, c0_n82_w72, c0_n82_w73, c0_n82_w74, c0_n82_w75, c0_n83_w1, c0_n83_w2, c0_n83_w3, c0_n83_w4, c0_n83_w5, c0_n83_w6, c0_n83_w7, c0_n83_w8, c0_n83_w9, c0_n83_w10, c0_n83_w11, c0_n83_w12, c0_n83_w13, c0_n83_w14, c0_n83_w15, c0_n83_w16, c0_n83_w17, c0_n83_w18, c0_n83_w19, c0_n83_w20, c0_n83_w21, c0_n83_w22, c0_n83_w23, c0_n83_w24, c0_n83_w25, c0_n83_w26, c0_n83_w27, c0_n83_w28, c0_n83_w29, c0_n83_w30, c0_n83_w31, c0_n83_w32, c0_n83_w33, c0_n83_w34, c0_n83_w35, c0_n83_w36, c0_n83_w37, c0_n83_w38, c0_n83_w39, c0_n83_w40, c0_n83_w41, c0_n83_w42, c0_n83_w43, c0_n83_w44, c0_n83_w45, c0_n83_w46, c0_n83_w47, c0_n83_w48, c0_n83_w49, c0_n83_w50, c0_n83_w51, c0_n83_w52, c0_n83_w53, c0_n83_w54, c0_n83_w55, c0_n83_w56, c0_n83_w57, c0_n83_w58, c0_n83_w59, c0_n83_w60, c0_n83_w61, c0_n83_w62, c0_n83_w63, c0_n83_w64, c0_n83_w65, c0_n83_w66, c0_n83_w67, c0_n83_w68, c0_n83_w69, c0_n83_w70, c0_n83_w71, c0_n83_w72, c0_n83_w73, c0_n83_w74, c0_n83_w75, c0_n84_w1, c0_n84_w2, c0_n84_w3, c0_n84_w4, c0_n84_w5, c0_n84_w6, c0_n84_w7, c0_n84_w8, c0_n84_w9, c0_n84_w10, c0_n84_w11, c0_n84_w12, c0_n84_w13, c0_n84_w14, c0_n84_w15, c0_n84_w16, c0_n84_w17, c0_n84_w18, c0_n84_w19, c0_n84_w20, c0_n84_w21, c0_n84_w22, c0_n84_w23, c0_n84_w24, c0_n84_w25, c0_n84_w26, c0_n84_w27, c0_n84_w28, c0_n84_w29, c0_n84_w30, c0_n84_w31, c0_n84_w32, c0_n84_w33, c0_n84_w34, c0_n84_w35, c0_n84_w36, c0_n84_w37, c0_n84_w38, c0_n84_w39, c0_n84_w40, c0_n84_w41, c0_n84_w42, c0_n84_w43, c0_n84_w44, c0_n84_w45, c0_n84_w46, c0_n84_w47, c0_n84_w48, c0_n84_w49, c0_n84_w50, c0_n84_w51, c0_n84_w52, c0_n84_w53, c0_n84_w54, c0_n84_w55, c0_n84_w56, c0_n84_w57, c0_n84_w58, c0_n84_w59, c0_n84_w60, c0_n84_w61, c0_n84_w62, c0_n84_w63, c0_n84_w64, c0_n84_w65, c0_n84_w66, c0_n84_w67, c0_n84_w68, c0_n84_w69, c0_n84_w70, c0_n84_w71, c0_n84_w72, c0_n84_w73, c0_n84_w74, c0_n84_w75, c0_n85_w1, c0_n85_w2, c0_n85_w3, c0_n85_w4, c0_n85_w5, c0_n85_w6, c0_n85_w7, c0_n85_w8, c0_n85_w9, c0_n85_w10, c0_n85_w11, c0_n85_w12, c0_n85_w13, c0_n85_w14, c0_n85_w15, c0_n85_w16, c0_n85_w17, c0_n85_w18, c0_n85_w19, c0_n85_w20, c0_n85_w21, c0_n85_w22, c0_n85_w23, c0_n85_w24, c0_n85_w25, c0_n85_w26, c0_n85_w27, c0_n85_w28, c0_n85_w29, c0_n85_w30, c0_n85_w31, c0_n85_w32, c0_n85_w33, c0_n85_w34, c0_n85_w35, c0_n85_w36, c0_n85_w37, c0_n85_w38, c0_n85_w39, c0_n85_w40, c0_n85_w41, c0_n85_w42, c0_n85_w43, c0_n85_w44, c0_n85_w45, c0_n85_w46, c0_n85_w47, c0_n85_w48, c0_n85_w49, c0_n85_w50, c0_n85_w51, c0_n85_w52, c0_n85_w53, c0_n85_w54, c0_n85_w55, c0_n85_w56, c0_n85_w57, c0_n85_w58, c0_n85_w59, c0_n85_w60, c0_n85_w61, c0_n85_w62, c0_n85_w63, c0_n85_w64, c0_n85_w65, c0_n85_w66, c0_n85_w67, c0_n85_w68, c0_n85_w69, c0_n85_w70, c0_n85_w71, c0_n85_w72, c0_n85_w73, c0_n85_w74, c0_n85_w75, c0_n86_w1, c0_n86_w2, c0_n86_w3, c0_n86_w4, c0_n86_w5, c0_n86_w6, c0_n86_w7, c0_n86_w8, c0_n86_w9, c0_n86_w10, c0_n86_w11, c0_n86_w12, c0_n86_w13, c0_n86_w14, c0_n86_w15, c0_n86_w16, c0_n86_w17, c0_n86_w18, c0_n86_w19, c0_n86_w20, c0_n86_w21, c0_n86_w22, c0_n86_w23, c0_n86_w24, c0_n86_w25, c0_n86_w26, c0_n86_w27, c0_n86_w28, c0_n86_w29, c0_n86_w30, c0_n86_w31, c0_n86_w32, c0_n86_w33, c0_n86_w34, c0_n86_w35, c0_n86_w36, c0_n86_w37, c0_n86_w38, c0_n86_w39, c0_n86_w40, c0_n86_w41, c0_n86_w42, c0_n86_w43, c0_n86_w44, c0_n86_w45, c0_n86_w46, c0_n86_w47, c0_n86_w48, c0_n86_w49, c0_n86_w50, c0_n86_w51, c0_n86_w52, c0_n86_w53, c0_n86_w54, c0_n86_w55, c0_n86_w56, c0_n86_w57, c0_n86_w58, c0_n86_w59, c0_n86_w60, c0_n86_w61, c0_n86_w62, c0_n86_w63, c0_n86_w64, c0_n86_w65, c0_n86_w66, c0_n86_w67, c0_n86_w68, c0_n86_w69, c0_n86_w70, c0_n86_w71, c0_n86_w72, c0_n86_w73, c0_n86_w74, c0_n86_w75, c0_n87_w1, c0_n87_w2, c0_n87_w3, c0_n87_w4, c0_n87_w5, c0_n87_w6, c0_n87_w7, c0_n87_w8, c0_n87_w9, c0_n87_w10, c0_n87_w11, c0_n87_w12, c0_n87_w13, c0_n87_w14, c0_n87_w15, c0_n87_w16, c0_n87_w17, c0_n87_w18, c0_n87_w19, c0_n87_w20, c0_n87_w21, c0_n87_w22, c0_n87_w23, c0_n87_w24, c0_n87_w25, c0_n87_w26, c0_n87_w27, c0_n87_w28, c0_n87_w29, c0_n87_w30, c0_n87_w31, c0_n87_w32, c0_n87_w33, c0_n87_w34, c0_n87_w35, c0_n87_w36, c0_n87_w37, c0_n87_w38, c0_n87_w39, c0_n87_w40, c0_n87_w41, c0_n87_w42, c0_n87_w43, c0_n87_w44, c0_n87_w45, c0_n87_w46, c0_n87_w47, c0_n87_w48, c0_n87_w49, c0_n87_w50, c0_n87_w51, c0_n87_w52, c0_n87_w53, c0_n87_w54, c0_n87_w55, c0_n87_w56, c0_n87_w57, c0_n87_w58, c0_n87_w59, c0_n87_w60, c0_n87_w61, c0_n87_w62, c0_n87_w63, c0_n87_w64, c0_n87_w65, c0_n87_w66, c0_n87_w67, c0_n87_w68, c0_n87_w69, c0_n87_w70, c0_n87_w71, c0_n87_w72, c0_n87_w73, c0_n87_w74, c0_n87_w75, c0_n88_w1, c0_n88_w2, c0_n88_w3, c0_n88_w4, c0_n88_w5, c0_n88_w6, c0_n88_w7, c0_n88_w8, c0_n88_w9, c0_n88_w10, c0_n88_w11, c0_n88_w12, c0_n88_w13, c0_n88_w14, c0_n88_w15, c0_n88_w16, c0_n88_w17, c0_n88_w18, c0_n88_w19, c0_n88_w20, c0_n88_w21, c0_n88_w22, c0_n88_w23, c0_n88_w24, c0_n88_w25, c0_n88_w26, c0_n88_w27, c0_n88_w28, c0_n88_w29, c0_n88_w30, c0_n88_w31, c0_n88_w32, c0_n88_w33, c0_n88_w34, c0_n88_w35, c0_n88_w36, c0_n88_w37, c0_n88_w38, c0_n88_w39, c0_n88_w40, c0_n88_w41, c0_n88_w42, c0_n88_w43, c0_n88_w44, c0_n88_w45, c0_n88_w46, c0_n88_w47, c0_n88_w48, c0_n88_w49, c0_n88_w50, c0_n88_w51, c0_n88_w52, c0_n88_w53, c0_n88_w54, c0_n88_w55, c0_n88_w56, c0_n88_w57, c0_n88_w58, c0_n88_w59, c0_n88_w60, c0_n88_w61, c0_n88_w62, c0_n88_w63, c0_n88_w64, c0_n88_w65, c0_n88_w66, c0_n88_w67, c0_n88_w68, c0_n88_w69, c0_n88_w70, c0_n88_w71, c0_n88_w72, c0_n88_w73, c0_n88_w74, c0_n88_w75, c0_n89_w1, c0_n89_w2, c0_n89_w3, c0_n89_w4, c0_n89_w5, c0_n89_w6, c0_n89_w7, c0_n89_w8, c0_n89_w9, c0_n89_w10, c0_n89_w11, c0_n89_w12, c0_n89_w13, c0_n89_w14, c0_n89_w15, c0_n89_w16, c0_n89_w17, c0_n89_w18, c0_n89_w19, c0_n89_w20, c0_n89_w21, c0_n89_w22, c0_n89_w23, c0_n89_w24, c0_n89_w25, c0_n89_w26, c0_n89_w27, c0_n89_w28, c0_n89_w29, c0_n89_w30, c0_n89_w31, c0_n89_w32, c0_n89_w33, c0_n89_w34, c0_n89_w35, c0_n89_w36, c0_n89_w37, c0_n89_w38, c0_n89_w39, c0_n89_w40, c0_n89_w41, c0_n89_w42, c0_n89_w43, c0_n89_w44, c0_n89_w45, c0_n89_w46, c0_n89_w47, c0_n89_w48, c0_n89_w49, c0_n89_w50, c0_n89_w51, c0_n89_w52, c0_n89_w53, c0_n89_w54, c0_n89_w55, c0_n89_w56, c0_n89_w57, c0_n89_w58, c0_n89_w59, c0_n89_w60, c0_n89_w61, c0_n89_w62, c0_n89_w63, c0_n89_w64, c0_n89_w65, c0_n89_w66, c0_n89_w67, c0_n89_w68, c0_n89_w69, c0_n89_w70, c0_n89_w71, c0_n89_w72, c0_n89_w73, c0_n89_w74, c0_n89_w75, c0_n90_w1, c0_n90_w2, c0_n90_w3, c0_n90_w4, c0_n90_w5, c0_n90_w6, c0_n90_w7, c0_n90_w8, c0_n90_w9, c0_n90_w10, c0_n90_w11, c0_n90_w12, c0_n90_w13, c0_n90_w14, c0_n90_w15, c0_n90_w16, c0_n90_w17, c0_n90_w18, c0_n90_w19, c0_n90_w20, c0_n90_w21, c0_n90_w22, c0_n90_w23, c0_n90_w24, c0_n90_w25, c0_n90_w26, c0_n90_w27, c0_n90_w28, c0_n90_w29, c0_n90_w30, c0_n90_w31, c0_n90_w32, c0_n90_w33, c0_n90_w34, c0_n90_w35, c0_n90_w36, c0_n90_w37, c0_n90_w38, c0_n90_w39, c0_n90_w40, c0_n90_w41, c0_n90_w42, c0_n90_w43, c0_n90_w44, c0_n90_w45, c0_n90_w46, c0_n90_w47, c0_n90_w48, c0_n90_w49, c0_n90_w50, c0_n90_w51, c0_n90_w52, c0_n90_w53, c0_n90_w54, c0_n90_w55, c0_n90_w56, c0_n90_w57, c0_n90_w58, c0_n90_w59, c0_n90_w60, c0_n90_w61, c0_n90_w62, c0_n90_w63, c0_n90_w64, c0_n90_w65, c0_n90_w66, c0_n90_w67, c0_n90_w68, c0_n90_w69, c0_n90_w70, c0_n90_w71, c0_n90_w72, c0_n90_w73, c0_n90_w74, c0_n90_w75, c0_n91_w1, c0_n91_w2, c0_n91_w3, c0_n91_w4, c0_n91_w5, c0_n91_w6, c0_n91_w7, c0_n91_w8, c0_n91_w9, c0_n91_w10, c0_n91_w11, c0_n91_w12, c0_n91_w13, c0_n91_w14, c0_n91_w15, c0_n91_w16, c0_n91_w17, c0_n91_w18, c0_n91_w19, c0_n91_w20, c0_n91_w21, c0_n91_w22, c0_n91_w23, c0_n91_w24, c0_n91_w25, c0_n91_w26, c0_n91_w27, c0_n91_w28, c0_n91_w29, c0_n91_w30, c0_n91_w31, c0_n91_w32, c0_n91_w33, c0_n91_w34, c0_n91_w35, c0_n91_w36, c0_n91_w37, c0_n91_w38, c0_n91_w39, c0_n91_w40, c0_n91_w41, c0_n91_w42, c0_n91_w43, c0_n91_w44, c0_n91_w45, c0_n91_w46, c0_n91_w47, c0_n91_w48, c0_n91_w49, c0_n91_w50, c0_n91_w51, c0_n91_w52, c0_n91_w53, c0_n91_w54, c0_n91_w55, c0_n91_w56, c0_n91_w57, c0_n91_w58, c0_n91_w59, c0_n91_w60, c0_n91_w61, c0_n91_w62, c0_n91_w63, c0_n91_w64, c0_n91_w65, c0_n91_w66, c0_n91_w67, c0_n91_w68, c0_n91_w69, c0_n91_w70, c0_n91_w71, c0_n91_w72, c0_n91_w73, c0_n91_w74, c0_n91_w75, c0_n92_w1, c0_n92_w2, c0_n92_w3, c0_n92_w4, c0_n92_w5, c0_n92_w6, c0_n92_w7, c0_n92_w8, c0_n92_w9, c0_n92_w10, c0_n92_w11, c0_n92_w12, c0_n92_w13, c0_n92_w14, c0_n92_w15, c0_n92_w16, c0_n92_w17, c0_n92_w18, c0_n92_w19, c0_n92_w20, c0_n92_w21, c0_n92_w22, c0_n92_w23, c0_n92_w24, c0_n92_w25, c0_n92_w26, c0_n92_w27, c0_n92_w28, c0_n92_w29, c0_n92_w30, c0_n92_w31, c0_n92_w32, c0_n92_w33, c0_n92_w34, c0_n92_w35, c0_n92_w36, c0_n92_w37, c0_n92_w38, c0_n92_w39, c0_n92_w40, c0_n92_w41, c0_n92_w42, c0_n92_w43, c0_n92_w44, c0_n92_w45, c0_n92_w46, c0_n92_w47, c0_n92_w48, c0_n92_w49, c0_n92_w50, c0_n92_w51, c0_n92_w52, c0_n92_w53, c0_n92_w54, c0_n92_w55, c0_n92_w56, c0_n92_w57, c0_n92_w58, c0_n92_w59, c0_n92_w60, c0_n92_w61, c0_n92_w62, c0_n92_w63, c0_n92_w64, c0_n92_w65, c0_n92_w66, c0_n92_w67, c0_n92_w68, c0_n92_w69, c0_n92_w70, c0_n92_w71, c0_n92_w72, c0_n92_w73, c0_n92_w74, c0_n92_w75, c0_n93_w1, c0_n93_w2, c0_n93_w3, c0_n93_w4, c0_n93_w5, c0_n93_w6, c0_n93_w7, c0_n93_w8, c0_n93_w9, c0_n93_w10, c0_n93_w11, c0_n93_w12, c0_n93_w13, c0_n93_w14, c0_n93_w15, c0_n93_w16, c0_n93_w17, c0_n93_w18, c0_n93_w19, c0_n93_w20, c0_n93_w21, c0_n93_w22, c0_n93_w23, c0_n93_w24, c0_n93_w25, c0_n93_w26, c0_n93_w27, c0_n93_w28, c0_n93_w29, c0_n93_w30, c0_n93_w31, c0_n93_w32, c0_n93_w33, c0_n93_w34, c0_n93_w35, c0_n93_w36, c0_n93_w37, c0_n93_w38, c0_n93_w39, c0_n93_w40, c0_n93_w41, c0_n93_w42, c0_n93_w43, c0_n93_w44, c0_n93_w45, c0_n93_w46, c0_n93_w47, c0_n93_w48, c0_n93_w49, c0_n93_w50, c0_n93_w51, c0_n93_w52, c0_n93_w53, c0_n93_w54, c0_n93_w55, c0_n93_w56, c0_n93_w57, c0_n93_w58, c0_n93_w59, c0_n93_w60, c0_n93_w61, c0_n93_w62, c0_n93_w63, c0_n93_w64, c0_n93_w65, c0_n93_w66, c0_n93_w67, c0_n93_w68, c0_n93_w69, c0_n93_w70, c0_n93_w71, c0_n93_w72, c0_n93_w73, c0_n93_w74, c0_n93_w75, c0_n94_w1, c0_n94_w2, c0_n94_w3, c0_n94_w4, c0_n94_w5, c0_n94_w6, c0_n94_w7, c0_n94_w8, c0_n94_w9, c0_n94_w10, c0_n94_w11, c0_n94_w12, c0_n94_w13, c0_n94_w14, c0_n94_w15, c0_n94_w16, c0_n94_w17, c0_n94_w18, c0_n94_w19, c0_n94_w20, c0_n94_w21, c0_n94_w22, c0_n94_w23, c0_n94_w24, c0_n94_w25, c0_n94_w26, c0_n94_w27, c0_n94_w28, c0_n94_w29, c0_n94_w30, c0_n94_w31, c0_n94_w32, c0_n94_w33, c0_n94_w34, c0_n94_w35, c0_n94_w36, c0_n94_w37, c0_n94_w38, c0_n94_w39, c0_n94_w40, c0_n94_w41, c0_n94_w42, c0_n94_w43, c0_n94_w44, c0_n94_w45, c0_n94_w46, c0_n94_w47, c0_n94_w48, c0_n94_w49, c0_n94_w50, c0_n94_w51, c0_n94_w52, c0_n94_w53, c0_n94_w54, c0_n94_w55, c0_n94_w56, c0_n94_w57, c0_n94_w58, c0_n94_w59, c0_n94_w60, c0_n94_w61, c0_n94_w62, c0_n94_w63, c0_n94_w64, c0_n94_w65, c0_n94_w66, c0_n94_w67, c0_n94_w68, c0_n94_w69, c0_n94_w70, c0_n94_w71, c0_n94_w72, c0_n94_w73, c0_n94_w74, c0_n94_w75, c0_n95_w1, c0_n95_w2, c0_n95_w3, c0_n95_w4, c0_n95_w5, c0_n95_w6, c0_n95_w7, c0_n95_w8, c0_n95_w9, c0_n95_w10, c0_n95_w11, c0_n95_w12, c0_n95_w13, c0_n95_w14, c0_n95_w15, c0_n95_w16, c0_n95_w17, c0_n95_w18, c0_n95_w19, c0_n95_w20, c0_n95_w21, c0_n95_w22, c0_n95_w23, c0_n95_w24, c0_n95_w25, c0_n95_w26, c0_n95_w27, c0_n95_w28, c0_n95_w29, c0_n95_w30, c0_n95_w31, c0_n95_w32, c0_n95_w33, c0_n95_w34, c0_n95_w35, c0_n95_w36, c0_n95_w37, c0_n95_w38, c0_n95_w39, c0_n95_w40, c0_n95_w41, c0_n95_w42, c0_n95_w43, c0_n95_w44, c0_n95_w45, c0_n95_w46, c0_n95_w47, c0_n95_w48, c0_n95_w49, c0_n95_w50, c0_n95_w51, c0_n95_w52, c0_n95_w53, c0_n95_w54, c0_n95_w55, c0_n95_w56, c0_n95_w57, c0_n95_w58, c0_n95_w59, c0_n95_w60, c0_n95_w61, c0_n95_w62, c0_n95_w63, c0_n95_w64, c0_n95_w65, c0_n95_w66, c0_n95_w67, c0_n95_w68, c0_n95_w69, c0_n95_w70, c0_n95_w71, c0_n95_w72, c0_n95_w73, c0_n95_w74, c0_n95_w75, c0_n96_w1, c0_n96_w2, c0_n96_w3, c0_n96_w4, c0_n96_w5, c0_n96_w6, c0_n96_w7, c0_n96_w8, c0_n96_w9, c0_n96_w10, c0_n96_w11, c0_n96_w12, c0_n96_w13, c0_n96_w14, c0_n96_w15, c0_n96_w16, c0_n96_w17, c0_n96_w18, c0_n96_w19, c0_n96_w20, c0_n96_w21, c0_n96_w22, c0_n96_w23, c0_n96_w24, c0_n96_w25, c0_n96_w26, c0_n96_w27, c0_n96_w28, c0_n96_w29, c0_n96_w30, c0_n96_w31, c0_n96_w32, c0_n96_w33, c0_n96_w34, c0_n96_w35, c0_n96_w36, c0_n96_w37, c0_n96_w38, c0_n96_w39, c0_n96_w40, c0_n96_w41, c0_n96_w42, c0_n96_w43, c0_n96_w44, c0_n96_w45, c0_n96_w46, c0_n96_w47, c0_n96_w48, c0_n96_w49, c0_n96_w50, c0_n96_w51, c0_n96_w52, c0_n96_w53, c0_n96_w54, c0_n96_w55, c0_n96_w56, c0_n96_w57, c0_n96_w58, c0_n96_w59, c0_n96_w60, c0_n96_w61, c0_n96_w62, c0_n96_w63, c0_n96_w64, c0_n96_w65, c0_n96_w66, c0_n96_w67, c0_n96_w68, c0_n96_w69, c0_n96_w70, c0_n96_w71, c0_n96_w72, c0_n96_w73, c0_n96_w74, c0_n96_w75, c0_n97_w1, c0_n97_w2, c0_n97_w3, c0_n97_w4, c0_n97_w5, c0_n97_w6, c0_n97_w7, c0_n97_w8, c0_n97_w9, c0_n97_w10, c0_n97_w11, c0_n97_w12, c0_n97_w13, c0_n97_w14, c0_n97_w15, c0_n97_w16, c0_n97_w17, c0_n97_w18, c0_n97_w19, c0_n97_w20, c0_n97_w21, c0_n97_w22, c0_n97_w23, c0_n97_w24, c0_n97_w25, c0_n97_w26, c0_n97_w27, c0_n97_w28, c0_n97_w29, c0_n97_w30, c0_n97_w31, c0_n97_w32, c0_n97_w33, c0_n97_w34, c0_n97_w35, c0_n97_w36, c0_n97_w37, c0_n97_w38, c0_n97_w39, c0_n97_w40, c0_n97_w41, c0_n97_w42, c0_n97_w43, c0_n97_w44, c0_n97_w45, c0_n97_w46, c0_n97_w47, c0_n97_w48, c0_n97_w49, c0_n97_w50, c0_n97_w51, c0_n97_w52, c0_n97_w53, c0_n97_w54, c0_n97_w55, c0_n97_w56, c0_n97_w57, c0_n97_w58, c0_n97_w59, c0_n97_w60, c0_n97_w61, c0_n97_w62, c0_n97_w63, c0_n97_w64, c0_n97_w65, c0_n97_w66, c0_n97_w67, c0_n97_w68, c0_n97_w69, c0_n97_w70, c0_n97_w71, c0_n97_w72, c0_n97_w73, c0_n97_w74, c0_n97_w75, c0_n98_w1, c0_n98_w2, c0_n98_w3, c0_n98_w4, c0_n98_w5, c0_n98_w6, c0_n98_w7, c0_n98_w8, c0_n98_w9, c0_n98_w10, c0_n98_w11, c0_n98_w12, c0_n98_w13, c0_n98_w14, c0_n98_w15, c0_n98_w16, c0_n98_w17, c0_n98_w18, c0_n98_w19, c0_n98_w20, c0_n98_w21, c0_n98_w22, c0_n98_w23, c0_n98_w24, c0_n98_w25, c0_n98_w26, c0_n98_w27, c0_n98_w28, c0_n98_w29, c0_n98_w30, c0_n98_w31, c0_n98_w32, c0_n98_w33, c0_n98_w34, c0_n98_w35, c0_n98_w36, c0_n98_w37, c0_n98_w38, c0_n98_w39, c0_n98_w40, c0_n98_w41, c0_n98_w42, c0_n98_w43, c0_n98_w44, c0_n98_w45, c0_n98_w46, c0_n98_w47, c0_n98_w48, c0_n98_w49, c0_n98_w50, c0_n98_w51, c0_n98_w52, c0_n98_w53, c0_n98_w54, c0_n98_w55, c0_n98_w56, c0_n98_w57, c0_n98_w58, c0_n98_w59, c0_n98_w60, c0_n98_w61, c0_n98_w62, c0_n98_w63, c0_n98_w64, c0_n98_w65, c0_n98_w66, c0_n98_w67, c0_n98_w68, c0_n98_w69, c0_n98_w70, c0_n98_w71, c0_n98_w72, c0_n98_w73, c0_n98_w74, c0_n98_w75, c0_n99_w1, c0_n99_w2, c0_n99_w3, c0_n99_w4, c0_n99_w5, c0_n99_w6, c0_n99_w7, c0_n99_w8, c0_n99_w9, c0_n99_w10, c0_n99_w11, c0_n99_w12, c0_n99_w13, c0_n99_w14, c0_n99_w15, c0_n99_w16, c0_n99_w17, c0_n99_w18, c0_n99_w19, c0_n99_w20, c0_n99_w21, c0_n99_w22, c0_n99_w23, c0_n99_w24, c0_n99_w25, c0_n99_w26, c0_n99_w27, c0_n99_w28, c0_n99_w29, c0_n99_w30, c0_n99_w31, c0_n99_w32, c0_n99_w33, c0_n99_w34, c0_n99_w35, c0_n99_w36, c0_n99_w37, c0_n99_w38, c0_n99_w39, c0_n99_w40, c0_n99_w41, c0_n99_w42, c0_n99_w43, c0_n99_w44, c0_n99_w45, c0_n99_w46, c0_n99_w47, c0_n99_w48, c0_n99_w49, c0_n99_w50, c0_n99_w51, c0_n99_w52, c0_n99_w53, c0_n99_w54, c0_n99_w55, c0_n99_w56, c0_n99_w57, c0_n99_w58, c0_n99_w59, c0_n99_w60, c0_n99_w61, c0_n99_w62, c0_n99_w63, c0_n99_w64, c0_n99_w65, c0_n99_w66, c0_n99_w67, c0_n99_w68, c0_n99_w69, c0_n99_w70, c0_n99_w71, c0_n99_w72, c0_n99_w73, c0_n99_w74, c0_n99_w75: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c0_n0_y, c0_n1_y, c0_n2_y, c0_n3_y, c0_n4_y, c0_n5_y, c0_n6_y, c0_n7_y, c0_n8_y, c0_n9_y, c0_n10_y, c0_n11_y, c0_n12_y, c0_n13_y, c0_n14_y, c0_n15_y, c0_n16_y, c0_n17_y, c0_n18_y, c0_n19_y, c0_n20_y, c0_n21_y, c0_n22_y, c0_n23_y, c0_n24_y, c0_n25_y, c0_n26_y, c0_n27_y, c0_n28_y, c0_n29_y, c0_n30_y, c0_n31_y, c0_n32_y, c0_n33_y, c0_n34_y, c0_n35_y, c0_n36_y, c0_n37_y, c0_n38_y, c0_n39_y, c0_n40_y, c0_n41_y, c0_n42_y, c0_n43_y, c0_n44_y, c0_n45_y, c0_n46_y, c0_n47_y, c0_n48_y, c0_n49_y, c0_n50_y, c0_n51_y, c0_n52_y, c0_n53_y, c0_n54_y, c0_n55_y, c0_n56_y, c0_n57_y, c0_n58_y, c0_n59_y, c0_n60_y, c0_n61_y, c0_n62_y, c0_n63_y, c0_n64_y, c0_n65_y, c0_n66_y, c0_n67_y, c0_n68_y, c0_n69_y, c0_n70_y, c0_n71_y, c0_n72_y, c0_n73_y, c0_n74_y, c0_n75_y, c0_n76_y, c0_n77_y, c0_n78_y, c0_n79_y, c0_n80_y, c0_n81_y, c0_n82_y, c0_n83_y, c0_n84_y, c0_n85_y, c0_n86_y, c0_n87_y, c0_n88_y, c0_n89_y, c0_n90_y, c0_n91_y, c0_n92_y, c0_n93_y, c0_n94_y, c0_n95_y, c0_n96_y, c0_n97_y, c0_n98_y, c0_n99_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada0_Leaky_ReLU_100neuron_8bits_75n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n0_w1, 
            w2=> c0_n0_w2, 
            w3=> c0_n0_w3, 
            w4=> c0_n0_w4, 
            w5=> c0_n0_w5, 
            w6=> c0_n0_w6, 
            w7=> c0_n0_w7, 
            w8=> c0_n0_w8, 
            w9=> c0_n0_w9, 
            w10=> c0_n0_w10, 
            w11=> c0_n0_w11, 
            w12=> c0_n0_w12, 
            w13=> c0_n0_w13, 
            w14=> c0_n0_w14, 
            w15=> c0_n0_w15, 
            w16=> c0_n0_w16, 
            w17=> c0_n0_w17, 
            w18=> c0_n0_w18, 
            w19=> c0_n0_w19, 
            w20=> c0_n0_w20, 
            w21=> c0_n0_w21, 
            w22=> c0_n0_w22, 
            w23=> c0_n0_w23, 
            w24=> c0_n0_w24, 
            w25=> c0_n0_w25, 
            w26=> c0_n0_w26, 
            w27=> c0_n0_w27, 
            w28=> c0_n0_w28, 
            w29=> c0_n0_w29, 
            w30=> c0_n0_w30, 
            w31=> c0_n0_w31, 
            w32=> c0_n0_w32, 
            w33=> c0_n0_w33, 
            w34=> c0_n0_w34, 
            w35=> c0_n0_w35, 
            w36=> c0_n0_w36, 
            w37=> c0_n0_w37, 
            w38=> c0_n0_w38, 
            w39=> c0_n0_w39, 
            w40=> c0_n0_w40, 
            w41=> c0_n0_w41, 
            w42=> c0_n0_w42, 
            w43=> c0_n0_w43, 
            w44=> c0_n0_w44, 
            w45=> c0_n0_w45, 
            w46=> c0_n0_w46, 
            w47=> c0_n0_w47, 
            w48=> c0_n0_w48, 
            w49=> c0_n0_w49, 
            w50=> c0_n0_w50, 
            w51=> c0_n0_w51, 
            w52=> c0_n0_w52, 
            w53=> c0_n0_w53, 
            w54=> c0_n0_w54, 
            w55=> c0_n0_w55, 
            w56=> c0_n0_w56, 
            w57=> c0_n0_w57, 
            w58=> c0_n0_w58, 
            w59=> c0_n0_w59, 
            w60=> c0_n0_w60, 
            w61=> c0_n0_w61, 
            w62=> c0_n0_w62, 
            w63=> c0_n0_w63, 
            w64=> c0_n0_w64, 
            w65=> c0_n0_w65, 
            w66=> c0_n0_w66, 
            w67=> c0_n0_w67, 
            w68=> c0_n0_w68, 
            w69=> c0_n0_w69, 
            w70=> c0_n0_w70, 
            w71=> c0_n0_w71, 
            w72=> c0_n0_w72, 
            w73=> c0_n0_w73, 
            w74=> c0_n0_w74, 
            w75=> c0_n0_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n1_w1, 
            w2=> c0_n1_w2, 
            w3=> c0_n1_w3, 
            w4=> c0_n1_w4, 
            w5=> c0_n1_w5, 
            w6=> c0_n1_w6, 
            w7=> c0_n1_w7, 
            w8=> c0_n1_w8, 
            w9=> c0_n1_w9, 
            w10=> c0_n1_w10, 
            w11=> c0_n1_w11, 
            w12=> c0_n1_w12, 
            w13=> c0_n1_w13, 
            w14=> c0_n1_w14, 
            w15=> c0_n1_w15, 
            w16=> c0_n1_w16, 
            w17=> c0_n1_w17, 
            w18=> c0_n1_w18, 
            w19=> c0_n1_w19, 
            w20=> c0_n1_w20, 
            w21=> c0_n1_w21, 
            w22=> c0_n1_w22, 
            w23=> c0_n1_w23, 
            w24=> c0_n1_w24, 
            w25=> c0_n1_w25, 
            w26=> c0_n1_w26, 
            w27=> c0_n1_w27, 
            w28=> c0_n1_w28, 
            w29=> c0_n1_w29, 
            w30=> c0_n1_w30, 
            w31=> c0_n1_w31, 
            w32=> c0_n1_w32, 
            w33=> c0_n1_w33, 
            w34=> c0_n1_w34, 
            w35=> c0_n1_w35, 
            w36=> c0_n1_w36, 
            w37=> c0_n1_w37, 
            w38=> c0_n1_w38, 
            w39=> c0_n1_w39, 
            w40=> c0_n1_w40, 
            w41=> c0_n1_w41, 
            w42=> c0_n1_w42, 
            w43=> c0_n1_w43, 
            w44=> c0_n1_w44, 
            w45=> c0_n1_w45, 
            w46=> c0_n1_w46, 
            w47=> c0_n1_w47, 
            w48=> c0_n1_w48, 
            w49=> c0_n1_w49, 
            w50=> c0_n1_w50, 
            w51=> c0_n1_w51, 
            w52=> c0_n1_w52, 
            w53=> c0_n1_w53, 
            w54=> c0_n1_w54, 
            w55=> c0_n1_w55, 
            w56=> c0_n1_w56, 
            w57=> c0_n1_w57, 
            w58=> c0_n1_w58, 
            w59=> c0_n1_w59, 
            w60=> c0_n1_w60, 
            w61=> c0_n1_w61, 
            w62=> c0_n1_w62, 
            w63=> c0_n1_w63, 
            w64=> c0_n1_w64, 
            w65=> c0_n1_w65, 
            w66=> c0_n1_w66, 
            w67=> c0_n1_w67, 
            w68=> c0_n1_w68, 
            w69=> c0_n1_w69, 
            w70=> c0_n1_w70, 
            w71=> c0_n1_w71, 
            w72=> c0_n1_w72, 
            w73=> c0_n1_w73, 
            w74=> c0_n1_w74, 
            w75=> c0_n1_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n2_w1, 
            w2=> c0_n2_w2, 
            w3=> c0_n2_w3, 
            w4=> c0_n2_w4, 
            w5=> c0_n2_w5, 
            w6=> c0_n2_w6, 
            w7=> c0_n2_w7, 
            w8=> c0_n2_w8, 
            w9=> c0_n2_w9, 
            w10=> c0_n2_w10, 
            w11=> c0_n2_w11, 
            w12=> c0_n2_w12, 
            w13=> c0_n2_w13, 
            w14=> c0_n2_w14, 
            w15=> c0_n2_w15, 
            w16=> c0_n2_w16, 
            w17=> c0_n2_w17, 
            w18=> c0_n2_w18, 
            w19=> c0_n2_w19, 
            w20=> c0_n2_w20, 
            w21=> c0_n2_w21, 
            w22=> c0_n2_w22, 
            w23=> c0_n2_w23, 
            w24=> c0_n2_w24, 
            w25=> c0_n2_w25, 
            w26=> c0_n2_w26, 
            w27=> c0_n2_w27, 
            w28=> c0_n2_w28, 
            w29=> c0_n2_w29, 
            w30=> c0_n2_w30, 
            w31=> c0_n2_w31, 
            w32=> c0_n2_w32, 
            w33=> c0_n2_w33, 
            w34=> c0_n2_w34, 
            w35=> c0_n2_w35, 
            w36=> c0_n2_w36, 
            w37=> c0_n2_w37, 
            w38=> c0_n2_w38, 
            w39=> c0_n2_w39, 
            w40=> c0_n2_w40, 
            w41=> c0_n2_w41, 
            w42=> c0_n2_w42, 
            w43=> c0_n2_w43, 
            w44=> c0_n2_w44, 
            w45=> c0_n2_w45, 
            w46=> c0_n2_w46, 
            w47=> c0_n2_w47, 
            w48=> c0_n2_w48, 
            w49=> c0_n2_w49, 
            w50=> c0_n2_w50, 
            w51=> c0_n2_w51, 
            w52=> c0_n2_w52, 
            w53=> c0_n2_w53, 
            w54=> c0_n2_w54, 
            w55=> c0_n2_w55, 
            w56=> c0_n2_w56, 
            w57=> c0_n2_w57, 
            w58=> c0_n2_w58, 
            w59=> c0_n2_w59, 
            w60=> c0_n2_w60, 
            w61=> c0_n2_w61, 
            w62=> c0_n2_w62, 
            w63=> c0_n2_w63, 
            w64=> c0_n2_w64, 
            w65=> c0_n2_w65, 
            w66=> c0_n2_w66, 
            w67=> c0_n2_w67, 
            w68=> c0_n2_w68, 
            w69=> c0_n2_w69, 
            w70=> c0_n2_w70, 
            w71=> c0_n2_w71, 
            w72=> c0_n2_w72, 
            w73=> c0_n2_w73, 
            w74=> c0_n2_w74, 
            w75=> c0_n2_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n3_w1, 
            w2=> c0_n3_w2, 
            w3=> c0_n3_w3, 
            w4=> c0_n3_w4, 
            w5=> c0_n3_w5, 
            w6=> c0_n3_w6, 
            w7=> c0_n3_w7, 
            w8=> c0_n3_w8, 
            w9=> c0_n3_w9, 
            w10=> c0_n3_w10, 
            w11=> c0_n3_w11, 
            w12=> c0_n3_w12, 
            w13=> c0_n3_w13, 
            w14=> c0_n3_w14, 
            w15=> c0_n3_w15, 
            w16=> c0_n3_w16, 
            w17=> c0_n3_w17, 
            w18=> c0_n3_w18, 
            w19=> c0_n3_w19, 
            w20=> c0_n3_w20, 
            w21=> c0_n3_w21, 
            w22=> c0_n3_w22, 
            w23=> c0_n3_w23, 
            w24=> c0_n3_w24, 
            w25=> c0_n3_w25, 
            w26=> c0_n3_w26, 
            w27=> c0_n3_w27, 
            w28=> c0_n3_w28, 
            w29=> c0_n3_w29, 
            w30=> c0_n3_w30, 
            w31=> c0_n3_w31, 
            w32=> c0_n3_w32, 
            w33=> c0_n3_w33, 
            w34=> c0_n3_w34, 
            w35=> c0_n3_w35, 
            w36=> c0_n3_w36, 
            w37=> c0_n3_w37, 
            w38=> c0_n3_w38, 
            w39=> c0_n3_w39, 
            w40=> c0_n3_w40, 
            w41=> c0_n3_w41, 
            w42=> c0_n3_w42, 
            w43=> c0_n3_w43, 
            w44=> c0_n3_w44, 
            w45=> c0_n3_w45, 
            w46=> c0_n3_w46, 
            w47=> c0_n3_w47, 
            w48=> c0_n3_w48, 
            w49=> c0_n3_w49, 
            w50=> c0_n3_w50, 
            w51=> c0_n3_w51, 
            w52=> c0_n3_w52, 
            w53=> c0_n3_w53, 
            w54=> c0_n3_w54, 
            w55=> c0_n3_w55, 
            w56=> c0_n3_w56, 
            w57=> c0_n3_w57, 
            w58=> c0_n3_w58, 
            w59=> c0_n3_w59, 
            w60=> c0_n3_w60, 
            w61=> c0_n3_w61, 
            w62=> c0_n3_w62, 
            w63=> c0_n3_w63, 
            w64=> c0_n3_w64, 
            w65=> c0_n3_w65, 
            w66=> c0_n3_w66, 
            w67=> c0_n3_w67, 
            w68=> c0_n3_w68, 
            w69=> c0_n3_w69, 
            w70=> c0_n3_w70, 
            w71=> c0_n3_w71, 
            w72=> c0_n3_w72, 
            w73=> c0_n3_w73, 
            w74=> c0_n3_w74, 
            w75=> c0_n3_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n4_w1, 
            w2=> c0_n4_w2, 
            w3=> c0_n4_w3, 
            w4=> c0_n4_w4, 
            w5=> c0_n4_w5, 
            w6=> c0_n4_w6, 
            w7=> c0_n4_w7, 
            w8=> c0_n4_w8, 
            w9=> c0_n4_w9, 
            w10=> c0_n4_w10, 
            w11=> c0_n4_w11, 
            w12=> c0_n4_w12, 
            w13=> c0_n4_w13, 
            w14=> c0_n4_w14, 
            w15=> c0_n4_w15, 
            w16=> c0_n4_w16, 
            w17=> c0_n4_w17, 
            w18=> c0_n4_w18, 
            w19=> c0_n4_w19, 
            w20=> c0_n4_w20, 
            w21=> c0_n4_w21, 
            w22=> c0_n4_w22, 
            w23=> c0_n4_w23, 
            w24=> c0_n4_w24, 
            w25=> c0_n4_w25, 
            w26=> c0_n4_w26, 
            w27=> c0_n4_w27, 
            w28=> c0_n4_w28, 
            w29=> c0_n4_w29, 
            w30=> c0_n4_w30, 
            w31=> c0_n4_w31, 
            w32=> c0_n4_w32, 
            w33=> c0_n4_w33, 
            w34=> c0_n4_w34, 
            w35=> c0_n4_w35, 
            w36=> c0_n4_w36, 
            w37=> c0_n4_w37, 
            w38=> c0_n4_w38, 
            w39=> c0_n4_w39, 
            w40=> c0_n4_w40, 
            w41=> c0_n4_w41, 
            w42=> c0_n4_w42, 
            w43=> c0_n4_w43, 
            w44=> c0_n4_w44, 
            w45=> c0_n4_w45, 
            w46=> c0_n4_w46, 
            w47=> c0_n4_w47, 
            w48=> c0_n4_w48, 
            w49=> c0_n4_w49, 
            w50=> c0_n4_w50, 
            w51=> c0_n4_w51, 
            w52=> c0_n4_w52, 
            w53=> c0_n4_w53, 
            w54=> c0_n4_w54, 
            w55=> c0_n4_w55, 
            w56=> c0_n4_w56, 
            w57=> c0_n4_w57, 
            w58=> c0_n4_w58, 
            w59=> c0_n4_w59, 
            w60=> c0_n4_w60, 
            w61=> c0_n4_w61, 
            w62=> c0_n4_w62, 
            w63=> c0_n4_w63, 
            w64=> c0_n4_w64, 
            w65=> c0_n4_w65, 
            w66=> c0_n4_w66, 
            w67=> c0_n4_w67, 
            w68=> c0_n4_w68, 
            w69=> c0_n4_w69, 
            w70=> c0_n4_w70, 
            w71=> c0_n4_w71, 
            w72=> c0_n4_w72, 
            w73=> c0_n4_w73, 
            w74=> c0_n4_w74, 
            w75=> c0_n4_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n5_w1, 
            w2=> c0_n5_w2, 
            w3=> c0_n5_w3, 
            w4=> c0_n5_w4, 
            w5=> c0_n5_w5, 
            w6=> c0_n5_w6, 
            w7=> c0_n5_w7, 
            w8=> c0_n5_w8, 
            w9=> c0_n5_w9, 
            w10=> c0_n5_w10, 
            w11=> c0_n5_w11, 
            w12=> c0_n5_w12, 
            w13=> c0_n5_w13, 
            w14=> c0_n5_w14, 
            w15=> c0_n5_w15, 
            w16=> c0_n5_w16, 
            w17=> c0_n5_w17, 
            w18=> c0_n5_w18, 
            w19=> c0_n5_w19, 
            w20=> c0_n5_w20, 
            w21=> c0_n5_w21, 
            w22=> c0_n5_w22, 
            w23=> c0_n5_w23, 
            w24=> c0_n5_w24, 
            w25=> c0_n5_w25, 
            w26=> c0_n5_w26, 
            w27=> c0_n5_w27, 
            w28=> c0_n5_w28, 
            w29=> c0_n5_w29, 
            w30=> c0_n5_w30, 
            w31=> c0_n5_w31, 
            w32=> c0_n5_w32, 
            w33=> c0_n5_w33, 
            w34=> c0_n5_w34, 
            w35=> c0_n5_w35, 
            w36=> c0_n5_w36, 
            w37=> c0_n5_w37, 
            w38=> c0_n5_w38, 
            w39=> c0_n5_w39, 
            w40=> c0_n5_w40, 
            w41=> c0_n5_w41, 
            w42=> c0_n5_w42, 
            w43=> c0_n5_w43, 
            w44=> c0_n5_w44, 
            w45=> c0_n5_w45, 
            w46=> c0_n5_w46, 
            w47=> c0_n5_w47, 
            w48=> c0_n5_w48, 
            w49=> c0_n5_w49, 
            w50=> c0_n5_w50, 
            w51=> c0_n5_w51, 
            w52=> c0_n5_w52, 
            w53=> c0_n5_w53, 
            w54=> c0_n5_w54, 
            w55=> c0_n5_w55, 
            w56=> c0_n5_w56, 
            w57=> c0_n5_w57, 
            w58=> c0_n5_w58, 
            w59=> c0_n5_w59, 
            w60=> c0_n5_w60, 
            w61=> c0_n5_w61, 
            w62=> c0_n5_w62, 
            w63=> c0_n5_w63, 
            w64=> c0_n5_w64, 
            w65=> c0_n5_w65, 
            w66=> c0_n5_w66, 
            w67=> c0_n5_w67, 
            w68=> c0_n5_w68, 
            w69=> c0_n5_w69, 
            w70=> c0_n5_w70, 
            w71=> c0_n5_w71, 
            w72=> c0_n5_w72, 
            w73=> c0_n5_w73, 
            w74=> c0_n5_w74, 
            w75=> c0_n5_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n6_w1, 
            w2=> c0_n6_w2, 
            w3=> c0_n6_w3, 
            w4=> c0_n6_w4, 
            w5=> c0_n6_w5, 
            w6=> c0_n6_w6, 
            w7=> c0_n6_w7, 
            w8=> c0_n6_w8, 
            w9=> c0_n6_w9, 
            w10=> c0_n6_w10, 
            w11=> c0_n6_w11, 
            w12=> c0_n6_w12, 
            w13=> c0_n6_w13, 
            w14=> c0_n6_w14, 
            w15=> c0_n6_w15, 
            w16=> c0_n6_w16, 
            w17=> c0_n6_w17, 
            w18=> c0_n6_w18, 
            w19=> c0_n6_w19, 
            w20=> c0_n6_w20, 
            w21=> c0_n6_w21, 
            w22=> c0_n6_w22, 
            w23=> c0_n6_w23, 
            w24=> c0_n6_w24, 
            w25=> c0_n6_w25, 
            w26=> c0_n6_w26, 
            w27=> c0_n6_w27, 
            w28=> c0_n6_w28, 
            w29=> c0_n6_w29, 
            w30=> c0_n6_w30, 
            w31=> c0_n6_w31, 
            w32=> c0_n6_w32, 
            w33=> c0_n6_w33, 
            w34=> c0_n6_w34, 
            w35=> c0_n6_w35, 
            w36=> c0_n6_w36, 
            w37=> c0_n6_w37, 
            w38=> c0_n6_w38, 
            w39=> c0_n6_w39, 
            w40=> c0_n6_w40, 
            w41=> c0_n6_w41, 
            w42=> c0_n6_w42, 
            w43=> c0_n6_w43, 
            w44=> c0_n6_w44, 
            w45=> c0_n6_w45, 
            w46=> c0_n6_w46, 
            w47=> c0_n6_w47, 
            w48=> c0_n6_w48, 
            w49=> c0_n6_w49, 
            w50=> c0_n6_w50, 
            w51=> c0_n6_w51, 
            w52=> c0_n6_w52, 
            w53=> c0_n6_w53, 
            w54=> c0_n6_w54, 
            w55=> c0_n6_w55, 
            w56=> c0_n6_w56, 
            w57=> c0_n6_w57, 
            w58=> c0_n6_w58, 
            w59=> c0_n6_w59, 
            w60=> c0_n6_w60, 
            w61=> c0_n6_w61, 
            w62=> c0_n6_w62, 
            w63=> c0_n6_w63, 
            w64=> c0_n6_w64, 
            w65=> c0_n6_w65, 
            w66=> c0_n6_w66, 
            w67=> c0_n6_w67, 
            w68=> c0_n6_w68, 
            w69=> c0_n6_w69, 
            w70=> c0_n6_w70, 
            w71=> c0_n6_w71, 
            w72=> c0_n6_w72, 
            w73=> c0_n6_w73, 
            w74=> c0_n6_w74, 
            w75=> c0_n6_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n7_w1, 
            w2=> c0_n7_w2, 
            w3=> c0_n7_w3, 
            w4=> c0_n7_w4, 
            w5=> c0_n7_w5, 
            w6=> c0_n7_w6, 
            w7=> c0_n7_w7, 
            w8=> c0_n7_w8, 
            w9=> c0_n7_w9, 
            w10=> c0_n7_w10, 
            w11=> c0_n7_w11, 
            w12=> c0_n7_w12, 
            w13=> c0_n7_w13, 
            w14=> c0_n7_w14, 
            w15=> c0_n7_w15, 
            w16=> c0_n7_w16, 
            w17=> c0_n7_w17, 
            w18=> c0_n7_w18, 
            w19=> c0_n7_w19, 
            w20=> c0_n7_w20, 
            w21=> c0_n7_w21, 
            w22=> c0_n7_w22, 
            w23=> c0_n7_w23, 
            w24=> c0_n7_w24, 
            w25=> c0_n7_w25, 
            w26=> c0_n7_w26, 
            w27=> c0_n7_w27, 
            w28=> c0_n7_w28, 
            w29=> c0_n7_w29, 
            w30=> c0_n7_w30, 
            w31=> c0_n7_w31, 
            w32=> c0_n7_w32, 
            w33=> c0_n7_w33, 
            w34=> c0_n7_w34, 
            w35=> c0_n7_w35, 
            w36=> c0_n7_w36, 
            w37=> c0_n7_w37, 
            w38=> c0_n7_w38, 
            w39=> c0_n7_w39, 
            w40=> c0_n7_w40, 
            w41=> c0_n7_w41, 
            w42=> c0_n7_w42, 
            w43=> c0_n7_w43, 
            w44=> c0_n7_w44, 
            w45=> c0_n7_w45, 
            w46=> c0_n7_w46, 
            w47=> c0_n7_w47, 
            w48=> c0_n7_w48, 
            w49=> c0_n7_w49, 
            w50=> c0_n7_w50, 
            w51=> c0_n7_w51, 
            w52=> c0_n7_w52, 
            w53=> c0_n7_w53, 
            w54=> c0_n7_w54, 
            w55=> c0_n7_w55, 
            w56=> c0_n7_w56, 
            w57=> c0_n7_w57, 
            w58=> c0_n7_w58, 
            w59=> c0_n7_w59, 
            w60=> c0_n7_w60, 
            w61=> c0_n7_w61, 
            w62=> c0_n7_w62, 
            w63=> c0_n7_w63, 
            w64=> c0_n7_w64, 
            w65=> c0_n7_w65, 
            w66=> c0_n7_w66, 
            w67=> c0_n7_w67, 
            w68=> c0_n7_w68, 
            w69=> c0_n7_w69, 
            w70=> c0_n7_w70, 
            w71=> c0_n7_w71, 
            w72=> c0_n7_w72, 
            w73=> c0_n7_w73, 
            w74=> c0_n7_w74, 
            w75=> c0_n7_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n8_w1, 
            w2=> c0_n8_w2, 
            w3=> c0_n8_w3, 
            w4=> c0_n8_w4, 
            w5=> c0_n8_w5, 
            w6=> c0_n8_w6, 
            w7=> c0_n8_w7, 
            w8=> c0_n8_w8, 
            w9=> c0_n8_w9, 
            w10=> c0_n8_w10, 
            w11=> c0_n8_w11, 
            w12=> c0_n8_w12, 
            w13=> c0_n8_w13, 
            w14=> c0_n8_w14, 
            w15=> c0_n8_w15, 
            w16=> c0_n8_w16, 
            w17=> c0_n8_w17, 
            w18=> c0_n8_w18, 
            w19=> c0_n8_w19, 
            w20=> c0_n8_w20, 
            w21=> c0_n8_w21, 
            w22=> c0_n8_w22, 
            w23=> c0_n8_w23, 
            w24=> c0_n8_w24, 
            w25=> c0_n8_w25, 
            w26=> c0_n8_w26, 
            w27=> c0_n8_w27, 
            w28=> c0_n8_w28, 
            w29=> c0_n8_w29, 
            w30=> c0_n8_w30, 
            w31=> c0_n8_w31, 
            w32=> c0_n8_w32, 
            w33=> c0_n8_w33, 
            w34=> c0_n8_w34, 
            w35=> c0_n8_w35, 
            w36=> c0_n8_w36, 
            w37=> c0_n8_w37, 
            w38=> c0_n8_w38, 
            w39=> c0_n8_w39, 
            w40=> c0_n8_w40, 
            w41=> c0_n8_w41, 
            w42=> c0_n8_w42, 
            w43=> c0_n8_w43, 
            w44=> c0_n8_w44, 
            w45=> c0_n8_w45, 
            w46=> c0_n8_w46, 
            w47=> c0_n8_w47, 
            w48=> c0_n8_w48, 
            w49=> c0_n8_w49, 
            w50=> c0_n8_w50, 
            w51=> c0_n8_w51, 
            w52=> c0_n8_w52, 
            w53=> c0_n8_w53, 
            w54=> c0_n8_w54, 
            w55=> c0_n8_w55, 
            w56=> c0_n8_w56, 
            w57=> c0_n8_w57, 
            w58=> c0_n8_w58, 
            w59=> c0_n8_w59, 
            w60=> c0_n8_w60, 
            w61=> c0_n8_w61, 
            w62=> c0_n8_w62, 
            w63=> c0_n8_w63, 
            w64=> c0_n8_w64, 
            w65=> c0_n8_w65, 
            w66=> c0_n8_w66, 
            w67=> c0_n8_w67, 
            w68=> c0_n8_w68, 
            w69=> c0_n8_w69, 
            w70=> c0_n8_w70, 
            w71=> c0_n8_w71, 
            w72=> c0_n8_w72, 
            w73=> c0_n8_w73, 
            w74=> c0_n8_w74, 
            w75=> c0_n8_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n9_w1, 
            w2=> c0_n9_w2, 
            w3=> c0_n9_w3, 
            w4=> c0_n9_w4, 
            w5=> c0_n9_w5, 
            w6=> c0_n9_w6, 
            w7=> c0_n9_w7, 
            w8=> c0_n9_w8, 
            w9=> c0_n9_w9, 
            w10=> c0_n9_w10, 
            w11=> c0_n9_w11, 
            w12=> c0_n9_w12, 
            w13=> c0_n9_w13, 
            w14=> c0_n9_w14, 
            w15=> c0_n9_w15, 
            w16=> c0_n9_w16, 
            w17=> c0_n9_w17, 
            w18=> c0_n9_w18, 
            w19=> c0_n9_w19, 
            w20=> c0_n9_w20, 
            w21=> c0_n9_w21, 
            w22=> c0_n9_w22, 
            w23=> c0_n9_w23, 
            w24=> c0_n9_w24, 
            w25=> c0_n9_w25, 
            w26=> c0_n9_w26, 
            w27=> c0_n9_w27, 
            w28=> c0_n9_w28, 
            w29=> c0_n9_w29, 
            w30=> c0_n9_w30, 
            w31=> c0_n9_w31, 
            w32=> c0_n9_w32, 
            w33=> c0_n9_w33, 
            w34=> c0_n9_w34, 
            w35=> c0_n9_w35, 
            w36=> c0_n9_w36, 
            w37=> c0_n9_w37, 
            w38=> c0_n9_w38, 
            w39=> c0_n9_w39, 
            w40=> c0_n9_w40, 
            w41=> c0_n9_w41, 
            w42=> c0_n9_w42, 
            w43=> c0_n9_w43, 
            w44=> c0_n9_w44, 
            w45=> c0_n9_w45, 
            w46=> c0_n9_w46, 
            w47=> c0_n9_w47, 
            w48=> c0_n9_w48, 
            w49=> c0_n9_w49, 
            w50=> c0_n9_w50, 
            w51=> c0_n9_w51, 
            w52=> c0_n9_w52, 
            w53=> c0_n9_w53, 
            w54=> c0_n9_w54, 
            w55=> c0_n9_w55, 
            w56=> c0_n9_w56, 
            w57=> c0_n9_w57, 
            w58=> c0_n9_w58, 
            w59=> c0_n9_w59, 
            w60=> c0_n9_w60, 
            w61=> c0_n9_w61, 
            w62=> c0_n9_w62, 
            w63=> c0_n9_w63, 
            w64=> c0_n9_w64, 
            w65=> c0_n9_w65, 
            w66=> c0_n9_w66, 
            w67=> c0_n9_w67, 
            w68=> c0_n9_w68, 
            w69=> c0_n9_w69, 
            w70=> c0_n9_w70, 
            w71=> c0_n9_w71, 
            w72=> c0_n9_w72, 
            w73=> c0_n9_w73, 
            w74=> c0_n9_w74, 
            w75=> c0_n9_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n9_y
   );           
            
neuron_inst_10: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n10_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n10_w1, 
            w2=> c0_n10_w2, 
            w3=> c0_n10_w3, 
            w4=> c0_n10_w4, 
            w5=> c0_n10_w5, 
            w6=> c0_n10_w6, 
            w7=> c0_n10_w7, 
            w8=> c0_n10_w8, 
            w9=> c0_n10_w9, 
            w10=> c0_n10_w10, 
            w11=> c0_n10_w11, 
            w12=> c0_n10_w12, 
            w13=> c0_n10_w13, 
            w14=> c0_n10_w14, 
            w15=> c0_n10_w15, 
            w16=> c0_n10_w16, 
            w17=> c0_n10_w17, 
            w18=> c0_n10_w18, 
            w19=> c0_n10_w19, 
            w20=> c0_n10_w20, 
            w21=> c0_n10_w21, 
            w22=> c0_n10_w22, 
            w23=> c0_n10_w23, 
            w24=> c0_n10_w24, 
            w25=> c0_n10_w25, 
            w26=> c0_n10_w26, 
            w27=> c0_n10_w27, 
            w28=> c0_n10_w28, 
            w29=> c0_n10_w29, 
            w30=> c0_n10_w30, 
            w31=> c0_n10_w31, 
            w32=> c0_n10_w32, 
            w33=> c0_n10_w33, 
            w34=> c0_n10_w34, 
            w35=> c0_n10_w35, 
            w36=> c0_n10_w36, 
            w37=> c0_n10_w37, 
            w38=> c0_n10_w38, 
            w39=> c0_n10_w39, 
            w40=> c0_n10_w40, 
            w41=> c0_n10_w41, 
            w42=> c0_n10_w42, 
            w43=> c0_n10_w43, 
            w44=> c0_n10_w44, 
            w45=> c0_n10_w45, 
            w46=> c0_n10_w46, 
            w47=> c0_n10_w47, 
            w48=> c0_n10_w48, 
            w49=> c0_n10_w49, 
            w50=> c0_n10_w50, 
            w51=> c0_n10_w51, 
            w52=> c0_n10_w52, 
            w53=> c0_n10_w53, 
            w54=> c0_n10_w54, 
            w55=> c0_n10_w55, 
            w56=> c0_n10_w56, 
            w57=> c0_n10_w57, 
            w58=> c0_n10_w58, 
            w59=> c0_n10_w59, 
            w60=> c0_n10_w60, 
            w61=> c0_n10_w61, 
            w62=> c0_n10_w62, 
            w63=> c0_n10_w63, 
            w64=> c0_n10_w64, 
            w65=> c0_n10_w65, 
            w66=> c0_n10_w66, 
            w67=> c0_n10_w67, 
            w68=> c0_n10_w68, 
            w69=> c0_n10_w69, 
            w70=> c0_n10_w70, 
            w71=> c0_n10_w71, 
            w72=> c0_n10_w72, 
            w73=> c0_n10_w73, 
            w74=> c0_n10_w74, 
            w75=> c0_n10_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n10_y
   );           
            
neuron_inst_11: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n11_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n11_w1, 
            w2=> c0_n11_w2, 
            w3=> c0_n11_w3, 
            w4=> c0_n11_w4, 
            w5=> c0_n11_w5, 
            w6=> c0_n11_w6, 
            w7=> c0_n11_w7, 
            w8=> c0_n11_w8, 
            w9=> c0_n11_w9, 
            w10=> c0_n11_w10, 
            w11=> c0_n11_w11, 
            w12=> c0_n11_w12, 
            w13=> c0_n11_w13, 
            w14=> c0_n11_w14, 
            w15=> c0_n11_w15, 
            w16=> c0_n11_w16, 
            w17=> c0_n11_w17, 
            w18=> c0_n11_w18, 
            w19=> c0_n11_w19, 
            w20=> c0_n11_w20, 
            w21=> c0_n11_w21, 
            w22=> c0_n11_w22, 
            w23=> c0_n11_w23, 
            w24=> c0_n11_w24, 
            w25=> c0_n11_w25, 
            w26=> c0_n11_w26, 
            w27=> c0_n11_w27, 
            w28=> c0_n11_w28, 
            w29=> c0_n11_w29, 
            w30=> c0_n11_w30, 
            w31=> c0_n11_w31, 
            w32=> c0_n11_w32, 
            w33=> c0_n11_w33, 
            w34=> c0_n11_w34, 
            w35=> c0_n11_w35, 
            w36=> c0_n11_w36, 
            w37=> c0_n11_w37, 
            w38=> c0_n11_w38, 
            w39=> c0_n11_w39, 
            w40=> c0_n11_w40, 
            w41=> c0_n11_w41, 
            w42=> c0_n11_w42, 
            w43=> c0_n11_w43, 
            w44=> c0_n11_w44, 
            w45=> c0_n11_w45, 
            w46=> c0_n11_w46, 
            w47=> c0_n11_w47, 
            w48=> c0_n11_w48, 
            w49=> c0_n11_w49, 
            w50=> c0_n11_w50, 
            w51=> c0_n11_w51, 
            w52=> c0_n11_w52, 
            w53=> c0_n11_w53, 
            w54=> c0_n11_w54, 
            w55=> c0_n11_w55, 
            w56=> c0_n11_w56, 
            w57=> c0_n11_w57, 
            w58=> c0_n11_w58, 
            w59=> c0_n11_w59, 
            w60=> c0_n11_w60, 
            w61=> c0_n11_w61, 
            w62=> c0_n11_w62, 
            w63=> c0_n11_w63, 
            w64=> c0_n11_w64, 
            w65=> c0_n11_w65, 
            w66=> c0_n11_w66, 
            w67=> c0_n11_w67, 
            w68=> c0_n11_w68, 
            w69=> c0_n11_w69, 
            w70=> c0_n11_w70, 
            w71=> c0_n11_w71, 
            w72=> c0_n11_w72, 
            w73=> c0_n11_w73, 
            w74=> c0_n11_w74, 
            w75=> c0_n11_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n11_y
   );           
            
neuron_inst_12: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n12_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n12_w1, 
            w2=> c0_n12_w2, 
            w3=> c0_n12_w3, 
            w4=> c0_n12_w4, 
            w5=> c0_n12_w5, 
            w6=> c0_n12_w6, 
            w7=> c0_n12_w7, 
            w8=> c0_n12_w8, 
            w9=> c0_n12_w9, 
            w10=> c0_n12_w10, 
            w11=> c0_n12_w11, 
            w12=> c0_n12_w12, 
            w13=> c0_n12_w13, 
            w14=> c0_n12_w14, 
            w15=> c0_n12_w15, 
            w16=> c0_n12_w16, 
            w17=> c0_n12_w17, 
            w18=> c0_n12_w18, 
            w19=> c0_n12_w19, 
            w20=> c0_n12_w20, 
            w21=> c0_n12_w21, 
            w22=> c0_n12_w22, 
            w23=> c0_n12_w23, 
            w24=> c0_n12_w24, 
            w25=> c0_n12_w25, 
            w26=> c0_n12_w26, 
            w27=> c0_n12_w27, 
            w28=> c0_n12_w28, 
            w29=> c0_n12_w29, 
            w30=> c0_n12_w30, 
            w31=> c0_n12_w31, 
            w32=> c0_n12_w32, 
            w33=> c0_n12_w33, 
            w34=> c0_n12_w34, 
            w35=> c0_n12_w35, 
            w36=> c0_n12_w36, 
            w37=> c0_n12_w37, 
            w38=> c0_n12_w38, 
            w39=> c0_n12_w39, 
            w40=> c0_n12_w40, 
            w41=> c0_n12_w41, 
            w42=> c0_n12_w42, 
            w43=> c0_n12_w43, 
            w44=> c0_n12_w44, 
            w45=> c0_n12_w45, 
            w46=> c0_n12_w46, 
            w47=> c0_n12_w47, 
            w48=> c0_n12_w48, 
            w49=> c0_n12_w49, 
            w50=> c0_n12_w50, 
            w51=> c0_n12_w51, 
            w52=> c0_n12_w52, 
            w53=> c0_n12_w53, 
            w54=> c0_n12_w54, 
            w55=> c0_n12_w55, 
            w56=> c0_n12_w56, 
            w57=> c0_n12_w57, 
            w58=> c0_n12_w58, 
            w59=> c0_n12_w59, 
            w60=> c0_n12_w60, 
            w61=> c0_n12_w61, 
            w62=> c0_n12_w62, 
            w63=> c0_n12_w63, 
            w64=> c0_n12_w64, 
            w65=> c0_n12_w65, 
            w66=> c0_n12_w66, 
            w67=> c0_n12_w67, 
            w68=> c0_n12_w68, 
            w69=> c0_n12_w69, 
            w70=> c0_n12_w70, 
            w71=> c0_n12_w71, 
            w72=> c0_n12_w72, 
            w73=> c0_n12_w73, 
            w74=> c0_n12_w74, 
            w75=> c0_n12_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n12_y
   );           
            
neuron_inst_13: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n13_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n13_w1, 
            w2=> c0_n13_w2, 
            w3=> c0_n13_w3, 
            w4=> c0_n13_w4, 
            w5=> c0_n13_w5, 
            w6=> c0_n13_w6, 
            w7=> c0_n13_w7, 
            w8=> c0_n13_w8, 
            w9=> c0_n13_w9, 
            w10=> c0_n13_w10, 
            w11=> c0_n13_w11, 
            w12=> c0_n13_w12, 
            w13=> c0_n13_w13, 
            w14=> c0_n13_w14, 
            w15=> c0_n13_w15, 
            w16=> c0_n13_w16, 
            w17=> c0_n13_w17, 
            w18=> c0_n13_w18, 
            w19=> c0_n13_w19, 
            w20=> c0_n13_w20, 
            w21=> c0_n13_w21, 
            w22=> c0_n13_w22, 
            w23=> c0_n13_w23, 
            w24=> c0_n13_w24, 
            w25=> c0_n13_w25, 
            w26=> c0_n13_w26, 
            w27=> c0_n13_w27, 
            w28=> c0_n13_w28, 
            w29=> c0_n13_w29, 
            w30=> c0_n13_w30, 
            w31=> c0_n13_w31, 
            w32=> c0_n13_w32, 
            w33=> c0_n13_w33, 
            w34=> c0_n13_w34, 
            w35=> c0_n13_w35, 
            w36=> c0_n13_w36, 
            w37=> c0_n13_w37, 
            w38=> c0_n13_w38, 
            w39=> c0_n13_w39, 
            w40=> c0_n13_w40, 
            w41=> c0_n13_w41, 
            w42=> c0_n13_w42, 
            w43=> c0_n13_w43, 
            w44=> c0_n13_w44, 
            w45=> c0_n13_w45, 
            w46=> c0_n13_w46, 
            w47=> c0_n13_w47, 
            w48=> c0_n13_w48, 
            w49=> c0_n13_w49, 
            w50=> c0_n13_w50, 
            w51=> c0_n13_w51, 
            w52=> c0_n13_w52, 
            w53=> c0_n13_w53, 
            w54=> c0_n13_w54, 
            w55=> c0_n13_w55, 
            w56=> c0_n13_w56, 
            w57=> c0_n13_w57, 
            w58=> c0_n13_w58, 
            w59=> c0_n13_w59, 
            w60=> c0_n13_w60, 
            w61=> c0_n13_w61, 
            w62=> c0_n13_w62, 
            w63=> c0_n13_w63, 
            w64=> c0_n13_w64, 
            w65=> c0_n13_w65, 
            w66=> c0_n13_w66, 
            w67=> c0_n13_w67, 
            w68=> c0_n13_w68, 
            w69=> c0_n13_w69, 
            w70=> c0_n13_w70, 
            w71=> c0_n13_w71, 
            w72=> c0_n13_w72, 
            w73=> c0_n13_w73, 
            w74=> c0_n13_w74, 
            w75=> c0_n13_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n13_y
   );           
            
neuron_inst_14: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n14_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n14_w1, 
            w2=> c0_n14_w2, 
            w3=> c0_n14_w3, 
            w4=> c0_n14_w4, 
            w5=> c0_n14_w5, 
            w6=> c0_n14_w6, 
            w7=> c0_n14_w7, 
            w8=> c0_n14_w8, 
            w9=> c0_n14_w9, 
            w10=> c0_n14_w10, 
            w11=> c0_n14_w11, 
            w12=> c0_n14_w12, 
            w13=> c0_n14_w13, 
            w14=> c0_n14_w14, 
            w15=> c0_n14_w15, 
            w16=> c0_n14_w16, 
            w17=> c0_n14_w17, 
            w18=> c0_n14_w18, 
            w19=> c0_n14_w19, 
            w20=> c0_n14_w20, 
            w21=> c0_n14_w21, 
            w22=> c0_n14_w22, 
            w23=> c0_n14_w23, 
            w24=> c0_n14_w24, 
            w25=> c0_n14_w25, 
            w26=> c0_n14_w26, 
            w27=> c0_n14_w27, 
            w28=> c0_n14_w28, 
            w29=> c0_n14_w29, 
            w30=> c0_n14_w30, 
            w31=> c0_n14_w31, 
            w32=> c0_n14_w32, 
            w33=> c0_n14_w33, 
            w34=> c0_n14_w34, 
            w35=> c0_n14_w35, 
            w36=> c0_n14_w36, 
            w37=> c0_n14_w37, 
            w38=> c0_n14_w38, 
            w39=> c0_n14_w39, 
            w40=> c0_n14_w40, 
            w41=> c0_n14_w41, 
            w42=> c0_n14_w42, 
            w43=> c0_n14_w43, 
            w44=> c0_n14_w44, 
            w45=> c0_n14_w45, 
            w46=> c0_n14_w46, 
            w47=> c0_n14_w47, 
            w48=> c0_n14_w48, 
            w49=> c0_n14_w49, 
            w50=> c0_n14_w50, 
            w51=> c0_n14_w51, 
            w52=> c0_n14_w52, 
            w53=> c0_n14_w53, 
            w54=> c0_n14_w54, 
            w55=> c0_n14_w55, 
            w56=> c0_n14_w56, 
            w57=> c0_n14_w57, 
            w58=> c0_n14_w58, 
            w59=> c0_n14_w59, 
            w60=> c0_n14_w60, 
            w61=> c0_n14_w61, 
            w62=> c0_n14_w62, 
            w63=> c0_n14_w63, 
            w64=> c0_n14_w64, 
            w65=> c0_n14_w65, 
            w66=> c0_n14_w66, 
            w67=> c0_n14_w67, 
            w68=> c0_n14_w68, 
            w69=> c0_n14_w69, 
            w70=> c0_n14_w70, 
            w71=> c0_n14_w71, 
            w72=> c0_n14_w72, 
            w73=> c0_n14_w73, 
            w74=> c0_n14_w74, 
            w75=> c0_n14_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n14_y
   );           
            
neuron_inst_15: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n15_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n15_w1, 
            w2=> c0_n15_w2, 
            w3=> c0_n15_w3, 
            w4=> c0_n15_w4, 
            w5=> c0_n15_w5, 
            w6=> c0_n15_w6, 
            w7=> c0_n15_w7, 
            w8=> c0_n15_w8, 
            w9=> c0_n15_w9, 
            w10=> c0_n15_w10, 
            w11=> c0_n15_w11, 
            w12=> c0_n15_w12, 
            w13=> c0_n15_w13, 
            w14=> c0_n15_w14, 
            w15=> c0_n15_w15, 
            w16=> c0_n15_w16, 
            w17=> c0_n15_w17, 
            w18=> c0_n15_w18, 
            w19=> c0_n15_w19, 
            w20=> c0_n15_w20, 
            w21=> c0_n15_w21, 
            w22=> c0_n15_w22, 
            w23=> c0_n15_w23, 
            w24=> c0_n15_w24, 
            w25=> c0_n15_w25, 
            w26=> c0_n15_w26, 
            w27=> c0_n15_w27, 
            w28=> c0_n15_w28, 
            w29=> c0_n15_w29, 
            w30=> c0_n15_w30, 
            w31=> c0_n15_w31, 
            w32=> c0_n15_w32, 
            w33=> c0_n15_w33, 
            w34=> c0_n15_w34, 
            w35=> c0_n15_w35, 
            w36=> c0_n15_w36, 
            w37=> c0_n15_w37, 
            w38=> c0_n15_w38, 
            w39=> c0_n15_w39, 
            w40=> c0_n15_w40, 
            w41=> c0_n15_w41, 
            w42=> c0_n15_w42, 
            w43=> c0_n15_w43, 
            w44=> c0_n15_w44, 
            w45=> c0_n15_w45, 
            w46=> c0_n15_w46, 
            w47=> c0_n15_w47, 
            w48=> c0_n15_w48, 
            w49=> c0_n15_w49, 
            w50=> c0_n15_w50, 
            w51=> c0_n15_w51, 
            w52=> c0_n15_w52, 
            w53=> c0_n15_w53, 
            w54=> c0_n15_w54, 
            w55=> c0_n15_w55, 
            w56=> c0_n15_w56, 
            w57=> c0_n15_w57, 
            w58=> c0_n15_w58, 
            w59=> c0_n15_w59, 
            w60=> c0_n15_w60, 
            w61=> c0_n15_w61, 
            w62=> c0_n15_w62, 
            w63=> c0_n15_w63, 
            w64=> c0_n15_w64, 
            w65=> c0_n15_w65, 
            w66=> c0_n15_w66, 
            w67=> c0_n15_w67, 
            w68=> c0_n15_w68, 
            w69=> c0_n15_w69, 
            w70=> c0_n15_w70, 
            w71=> c0_n15_w71, 
            w72=> c0_n15_w72, 
            w73=> c0_n15_w73, 
            w74=> c0_n15_w74, 
            w75=> c0_n15_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n15_y
   );           
            
neuron_inst_16: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n16_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n16_w1, 
            w2=> c0_n16_w2, 
            w3=> c0_n16_w3, 
            w4=> c0_n16_w4, 
            w5=> c0_n16_w5, 
            w6=> c0_n16_w6, 
            w7=> c0_n16_w7, 
            w8=> c0_n16_w8, 
            w9=> c0_n16_w9, 
            w10=> c0_n16_w10, 
            w11=> c0_n16_w11, 
            w12=> c0_n16_w12, 
            w13=> c0_n16_w13, 
            w14=> c0_n16_w14, 
            w15=> c0_n16_w15, 
            w16=> c0_n16_w16, 
            w17=> c0_n16_w17, 
            w18=> c0_n16_w18, 
            w19=> c0_n16_w19, 
            w20=> c0_n16_w20, 
            w21=> c0_n16_w21, 
            w22=> c0_n16_w22, 
            w23=> c0_n16_w23, 
            w24=> c0_n16_w24, 
            w25=> c0_n16_w25, 
            w26=> c0_n16_w26, 
            w27=> c0_n16_w27, 
            w28=> c0_n16_w28, 
            w29=> c0_n16_w29, 
            w30=> c0_n16_w30, 
            w31=> c0_n16_w31, 
            w32=> c0_n16_w32, 
            w33=> c0_n16_w33, 
            w34=> c0_n16_w34, 
            w35=> c0_n16_w35, 
            w36=> c0_n16_w36, 
            w37=> c0_n16_w37, 
            w38=> c0_n16_w38, 
            w39=> c0_n16_w39, 
            w40=> c0_n16_w40, 
            w41=> c0_n16_w41, 
            w42=> c0_n16_w42, 
            w43=> c0_n16_w43, 
            w44=> c0_n16_w44, 
            w45=> c0_n16_w45, 
            w46=> c0_n16_w46, 
            w47=> c0_n16_w47, 
            w48=> c0_n16_w48, 
            w49=> c0_n16_w49, 
            w50=> c0_n16_w50, 
            w51=> c0_n16_w51, 
            w52=> c0_n16_w52, 
            w53=> c0_n16_w53, 
            w54=> c0_n16_w54, 
            w55=> c0_n16_w55, 
            w56=> c0_n16_w56, 
            w57=> c0_n16_w57, 
            w58=> c0_n16_w58, 
            w59=> c0_n16_w59, 
            w60=> c0_n16_w60, 
            w61=> c0_n16_w61, 
            w62=> c0_n16_w62, 
            w63=> c0_n16_w63, 
            w64=> c0_n16_w64, 
            w65=> c0_n16_w65, 
            w66=> c0_n16_w66, 
            w67=> c0_n16_w67, 
            w68=> c0_n16_w68, 
            w69=> c0_n16_w69, 
            w70=> c0_n16_w70, 
            w71=> c0_n16_w71, 
            w72=> c0_n16_w72, 
            w73=> c0_n16_w73, 
            w74=> c0_n16_w74, 
            w75=> c0_n16_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n16_y
   );           
            
neuron_inst_17: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n17_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n17_w1, 
            w2=> c0_n17_w2, 
            w3=> c0_n17_w3, 
            w4=> c0_n17_w4, 
            w5=> c0_n17_w5, 
            w6=> c0_n17_w6, 
            w7=> c0_n17_w7, 
            w8=> c0_n17_w8, 
            w9=> c0_n17_w9, 
            w10=> c0_n17_w10, 
            w11=> c0_n17_w11, 
            w12=> c0_n17_w12, 
            w13=> c0_n17_w13, 
            w14=> c0_n17_w14, 
            w15=> c0_n17_w15, 
            w16=> c0_n17_w16, 
            w17=> c0_n17_w17, 
            w18=> c0_n17_w18, 
            w19=> c0_n17_w19, 
            w20=> c0_n17_w20, 
            w21=> c0_n17_w21, 
            w22=> c0_n17_w22, 
            w23=> c0_n17_w23, 
            w24=> c0_n17_w24, 
            w25=> c0_n17_w25, 
            w26=> c0_n17_w26, 
            w27=> c0_n17_w27, 
            w28=> c0_n17_w28, 
            w29=> c0_n17_w29, 
            w30=> c0_n17_w30, 
            w31=> c0_n17_w31, 
            w32=> c0_n17_w32, 
            w33=> c0_n17_w33, 
            w34=> c0_n17_w34, 
            w35=> c0_n17_w35, 
            w36=> c0_n17_w36, 
            w37=> c0_n17_w37, 
            w38=> c0_n17_w38, 
            w39=> c0_n17_w39, 
            w40=> c0_n17_w40, 
            w41=> c0_n17_w41, 
            w42=> c0_n17_w42, 
            w43=> c0_n17_w43, 
            w44=> c0_n17_w44, 
            w45=> c0_n17_w45, 
            w46=> c0_n17_w46, 
            w47=> c0_n17_w47, 
            w48=> c0_n17_w48, 
            w49=> c0_n17_w49, 
            w50=> c0_n17_w50, 
            w51=> c0_n17_w51, 
            w52=> c0_n17_w52, 
            w53=> c0_n17_w53, 
            w54=> c0_n17_w54, 
            w55=> c0_n17_w55, 
            w56=> c0_n17_w56, 
            w57=> c0_n17_w57, 
            w58=> c0_n17_w58, 
            w59=> c0_n17_w59, 
            w60=> c0_n17_w60, 
            w61=> c0_n17_w61, 
            w62=> c0_n17_w62, 
            w63=> c0_n17_w63, 
            w64=> c0_n17_w64, 
            w65=> c0_n17_w65, 
            w66=> c0_n17_w66, 
            w67=> c0_n17_w67, 
            w68=> c0_n17_w68, 
            w69=> c0_n17_w69, 
            w70=> c0_n17_w70, 
            w71=> c0_n17_w71, 
            w72=> c0_n17_w72, 
            w73=> c0_n17_w73, 
            w74=> c0_n17_w74, 
            w75=> c0_n17_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n17_y
   );           
            
neuron_inst_18: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n18_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n18_w1, 
            w2=> c0_n18_w2, 
            w3=> c0_n18_w3, 
            w4=> c0_n18_w4, 
            w5=> c0_n18_w5, 
            w6=> c0_n18_w6, 
            w7=> c0_n18_w7, 
            w8=> c0_n18_w8, 
            w9=> c0_n18_w9, 
            w10=> c0_n18_w10, 
            w11=> c0_n18_w11, 
            w12=> c0_n18_w12, 
            w13=> c0_n18_w13, 
            w14=> c0_n18_w14, 
            w15=> c0_n18_w15, 
            w16=> c0_n18_w16, 
            w17=> c0_n18_w17, 
            w18=> c0_n18_w18, 
            w19=> c0_n18_w19, 
            w20=> c0_n18_w20, 
            w21=> c0_n18_w21, 
            w22=> c0_n18_w22, 
            w23=> c0_n18_w23, 
            w24=> c0_n18_w24, 
            w25=> c0_n18_w25, 
            w26=> c0_n18_w26, 
            w27=> c0_n18_w27, 
            w28=> c0_n18_w28, 
            w29=> c0_n18_w29, 
            w30=> c0_n18_w30, 
            w31=> c0_n18_w31, 
            w32=> c0_n18_w32, 
            w33=> c0_n18_w33, 
            w34=> c0_n18_w34, 
            w35=> c0_n18_w35, 
            w36=> c0_n18_w36, 
            w37=> c0_n18_w37, 
            w38=> c0_n18_w38, 
            w39=> c0_n18_w39, 
            w40=> c0_n18_w40, 
            w41=> c0_n18_w41, 
            w42=> c0_n18_w42, 
            w43=> c0_n18_w43, 
            w44=> c0_n18_w44, 
            w45=> c0_n18_w45, 
            w46=> c0_n18_w46, 
            w47=> c0_n18_w47, 
            w48=> c0_n18_w48, 
            w49=> c0_n18_w49, 
            w50=> c0_n18_w50, 
            w51=> c0_n18_w51, 
            w52=> c0_n18_w52, 
            w53=> c0_n18_w53, 
            w54=> c0_n18_w54, 
            w55=> c0_n18_w55, 
            w56=> c0_n18_w56, 
            w57=> c0_n18_w57, 
            w58=> c0_n18_w58, 
            w59=> c0_n18_w59, 
            w60=> c0_n18_w60, 
            w61=> c0_n18_w61, 
            w62=> c0_n18_w62, 
            w63=> c0_n18_w63, 
            w64=> c0_n18_w64, 
            w65=> c0_n18_w65, 
            w66=> c0_n18_w66, 
            w67=> c0_n18_w67, 
            w68=> c0_n18_w68, 
            w69=> c0_n18_w69, 
            w70=> c0_n18_w70, 
            w71=> c0_n18_w71, 
            w72=> c0_n18_w72, 
            w73=> c0_n18_w73, 
            w74=> c0_n18_w74, 
            w75=> c0_n18_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n18_y
   );           
            
neuron_inst_19: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n19_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n19_w1, 
            w2=> c0_n19_w2, 
            w3=> c0_n19_w3, 
            w4=> c0_n19_w4, 
            w5=> c0_n19_w5, 
            w6=> c0_n19_w6, 
            w7=> c0_n19_w7, 
            w8=> c0_n19_w8, 
            w9=> c0_n19_w9, 
            w10=> c0_n19_w10, 
            w11=> c0_n19_w11, 
            w12=> c0_n19_w12, 
            w13=> c0_n19_w13, 
            w14=> c0_n19_w14, 
            w15=> c0_n19_w15, 
            w16=> c0_n19_w16, 
            w17=> c0_n19_w17, 
            w18=> c0_n19_w18, 
            w19=> c0_n19_w19, 
            w20=> c0_n19_w20, 
            w21=> c0_n19_w21, 
            w22=> c0_n19_w22, 
            w23=> c0_n19_w23, 
            w24=> c0_n19_w24, 
            w25=> c0_n19_w25, 
            w26=> c0_n19_w26, 
            w27=> c0_n19_w27, 
            w28=> c0_n19_w28, 
            w29=> c0_n19_w29, 
            w30=> c0_n19_w30, 
            w31=> c0_n19_w31, 
            w32=> c0_n19_w32, 
            w33=> c0_n19_w33, 
            w34=> c0_n19_w34, 
            w35=> c0_n19_w35, 
            w36=> c0_n19_w36, 
            w37=> c0_n19_w37, 
            w38=> c0_n19_w38, 
            w39=> c0_n19_w39, 
            w40=> c0_n19_w40, 
            w41=> c0_n19_w41, 
            w42=> c0_n19_w42, 
            w43=> c0_n19_w43, 
            w44=> c0_n19_w44, 
            w45=> c0_n19_w45, 
            w46=> c0_n19_w46, 
            w47=> c0_n19_w47, 
            w48=> c0_n19_w48, 
            w49=> c0_n19_w49, 
            w50=> c0_n19_w50, 
            w51=> c0_n19_w51, 
            w52=> c0_n19_w52, 
            w53=> c0_n19_w53, 
            w54=> c0_n19_w54, 
            w55=> c0_n19_w55, 
            w56=> c0_n19_w56, 
            w57=> c0_n19_w57, 
            w58=> c0_n19_w58, 
            w59=> c0_n19_w59, 
            w60=> c0_n19_w60, 
            w61=> c0_n19_w61, 
            w62=> c0_n19_w62, 
            w63=> c0_n19_w63, 
            w64=> c0_n19_w64, 
            w65=> c0_n19_w65, 
            w66=> c0_n19_w66, 
            w67=> c0_n19_w67, 
            w68=> c0_n19_w68, 
            w69=> c0_n19_w69, 
            w70=> c0_n19_w70, 
            w71=> c0_n19_w71, 
            w72=> c0_n19_w72, 
            w73=> c0_n19_w73, 
            w74=> c0_n19_w74, 
            w75=> c0_n19_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n19_y
   );           
            
neuron_inst_20: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n20_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n20_w1, 
            w2=> c0_n20_w2, 
            w3=> c0_n20_w3, 
            w4=> c0_n20_w4, 
            w5=> c0_n20_w5, 
            w6=> c0_n20_w6, 
            w7=> c0_n20_w7, 
            w8=> c0_n20_w8, 
            w9=> c0_n20_w9, 
            w10=> c0_n20_w10, 
            w11=> c0_n20_w11, 
            w12=> c0_n20_w12, 
            w13=> c0_n20_w13, 
            w14=> c0_n20_w14, 
            w15=> c0_n20_w15, 
            w16=> c0_n20_w16, 
            w17=> c0_n20_w17, 
            w18=> c0_n20_w18, 
            w19=> c0_n20_w19, 
            w20=> c0_n20_w20, 
            w21=> c0_n20_w21, 
            w22=> c0_n20_w22, 
            w23=> c0_n20_w23, 
            w24=> c0_n20_w24, 
            w25=> c0_n20_w25, 
            w26=> c0_n20_w26, 
            w27=> c0_n20_w27, 
            w28=> c0_n20_w28, 
            w29=> c0_n20_w29, 
            w30=> c0_n20_w30, 
            w31=> c0_n20_w31, 
            w32=> c0_n20_w32, 
            w33=> c0_n20_w33, 
            w34=> c0_n20_w34, 
            w35=> c0_n20_w35, 
            w36=> c0_n20_w36, 
            w37=> c0_n20_w37, 
            w38=> c0_n20_w38, 
            w39=> c0_n20_w39, 
            w40=> c0_n20_w40, 
            w41=> c0_n20_w41, 
            w42=> c0_n20_w42, 
            w43=> c0_n20_w43, 
            w44=> c0_n20_w44, 
            w45=> c0_n20_w45, 
            w46=> c0_n20_w46, 
            w47=> c0_n20_w47, 
            w48=> c0_n20_w48, 
            w49=> c0_n20_w49, 
            w50=> c0_n20_w50, 
            w51=> c0_n20_w51, 
            w52=> c0_n20_w52, 
            w53=> c0_n20_w53, 
            w54=> c0_n20_w54, 
            w55=> c0_n20_w55, 
            w56=> c0_n20_w56, 
            w57=> c0_n20_w57, 
            w58=> c0_n20_w58, 
            w59=> c0_n20_w59, 
            w60=> c0_n20_w60, 
            w61=> c0_n20_w61, 
            w62=> c0_n20_w62, 
            w63=> c0_n20_w63, 
            w64=> c0_n20_w64, 
            w65=> c0_n20_w65, 
            w66=> c0_n20_w66, 
            w67=> c0_n20_w67, 
            w68=> c0_n20_w68, 
            w69=> c0_n20_w69, 
            w70=> c0_n20_w70, 
            w71=> c0_n20_w71, 
            w72=> c0_n20_w72, 
            w73=> c0_n20_w73, 
            w74=> c0_n20_w74, 
            w75=> c0_n20_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n20_y
   );           
            
neuron_inst_21: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n21_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n21_w1, 
            w2=> c0_n21_w2, 
            w3=> c0_n21_w3, 
            w4=> c0_n21_w4, 
            w5=> c0_n21_w5, 
            w6=> c0_n21_w6, 
            w7=> c0_n21_w7, 
            w8=> c0_n21_w8, 
            w9=> c0_n21_w9, 
            w10=> c0_n21_w10, 
            w11=> c0_n21_w11, 
            w12=> c0_n21_w12, 
            w13=> c0_n21_w13, 
            w14=> c0_n21_w14, 
            w15=> c0_n21_w15, 
            w16=> c0_n21_w16, 
            w17=> c0_n21_w17, 
            w18=> c0_n21_w18, 
            w19=> c0_n21_w19, 
            w20=> c0_n21_w20, 
            w21=> c0_n21_w21, 
            w22=> c0_n21_w22, 
            w23=> c0_n21_w23, 
            w24=> c0_n21_w24, 
            w25=> c0_n21_w25, 
            w26=> c0_n21_w26, 
            w27=> c0_n21_w27, 
            w28=> c0_n21_w28, 
            w29=> c0_n21_w29, 
            w30=> c0_n21_w30, 
            w31=> c0_n21_w31, 
            w32=> c0_n21_w32, 
            w33=> c0_n21_w33, 
            w34=> c0_n21_w34, 
            w35=> c0_n21_w35, 
            w36=> c0_n21_w36, 
            w37=> c0_n21_w37, 
            w38=> c0_n21_w38, 
            w39=> c0_n21_w39, 
            w40=> c0_n21_w40, 
            w41=> c0_n21_w41, 
            w42=> c0_n21_w42, 
            w43=> c0_n21_w43, 
            w44=> c0_n21_w44, 
            w45=> c0_n21_w45, 
            w46=> c0_n21_w46, 
            w47=> c0_n21_w47, 
            w48=> c0_n21_w48, 
            w49=> c0_n21_w49, 
            w50=> c0_n21_w50, 
            w51=> c0_n21_w51, 
            w52=> c0_n21_w52, 
            w53=> c0_n21_w53, 
            w54=> c0_n21_w54, 
            w55=> c0_n21_w55, 
            w56=> c0_n21_w56, 
            w57=> c0_n21_w57, 
            w58=> c0_n21_w58, 
            w59=> c0_n21_w59, 
            w60=> c0_n21_w60, 
            w61=> c0_n21_w61, 
            w62=> c0_n21_w62, 
            w63=> c0_n21_w63, 
            w64=> c0_n21_w64, 
            w65=> c0_n21_w65, 
            w66=> c0_n21_w66, 
            w67=> c0_n21_w67, 
            w68=> c0_n21_w68, 
            w69=> c0_n21_w69, 
            w70=> c0_n21_w70, 
            w71=> c0_n21_w71, 
            w72=> c0_n21_w72, 
            w73=> c0_n21_w73, 
            w74=> c0_n21_w74, 
            w75=> c0_n21_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n21_y
   );           
            
neuron_inst_22: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n22_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n22_w1, 
            w2=> c0_n22_w2, 
            w3=> c0_n22_w3, 
            w4=> c0_n22_w4, 
            w5=> c0_n22_w5, 
            w6=> c0_n22_w6, 
            w7=> c0_n22_w7, 
            w8=> c0_n22_w8, 
            w9=> c0_n22_w9, 
            w10=> c0_n22_w10, 
            w11=> c0_n22_w11, 
            w12=> c0_n22_w12, 
            w13=> c0_n22_w13, 
            w14=> c0_n22_w14, 
            w15=> c0_n22_w15, 
            w16=> c0_n22_w16, 
            w17=> c0_n22_w17, 
            w18=> c0_n22_w18, 
            w19=> c0_n22_w19, 
            w20=> c0_n22_w20, 
            w21=> c0_n22_w21, 
            w22=> c0_n22_w22, 
            w23=> c0_n22_w23, 
            w24=> c0_n22_w24, 
            w25=> c0_n22_w25, 
            w26=> c0_n22_w26, 
            w27=> c0_n22_w27, 
            w28=> c0_n22_w28, 
            w29=> c0_n22_w29, 
            w30=> c0_n22_w30, 
            w31=> c0_n22_w31, 
            w32=> c0_n22_w32, 
            w33=> c0_n22_w33, 
            w34=> c0_n22_w34, 
            w35=> c0_n22_w35, 
            w36=> c0_n22_w36, 
            w37=> c0_n22_w37, 
            w38=> c0_n22_w38, 
            w39=> c0_n22_w39, 
            w40=> c0_n22_w40, 
            w41=> c0_n22_w41, 
            w42=> c0_n22_w42, 
            w43=> c0_n22_w43, 
            w44=> c0_n22_w44, 
            w45=> c0_n22_w45, 
            w46=> c0_n22_w46, 
            w47=> c0_n22_w47, 
            w48=> c0_n22_w48, 
            w49=> c0_n22_w49, 
            w50=> c0_n22_w50, 
            w51=> c0_n22_w51, 
            w52=> c0_n22_w52, 
            w53=> c0_n22_w53, 
            w54=> c0_n22_w54, 
            w55=> c0_n22_w55, 
            w56=> c0_n22_w56, 
            w57=> c0_n22_w57, 
            w58=> c0_n22_w58, 
            w59=> c0_n22_w59, 
            w60=> c0_n22_w60, 
            w61=> c0_n22_w61, 
            w62=> c0_n22_w62, 
            w63=> c0_n22_w63, 
            w64=> c0_n22_w64, 
            w65=> c0_n22_w65, 
            w66=> c0_n22_w66, 
            w67=> c0_n22_w67, 
            w68=> c0_n22_w68, 
            w69=> c0_n22_w69, 
            w70=> c0_n22_w70, 
            w71=> c0_n22_w71, 
            w72=> c0_n22_w72, 
            w73=> c0_n22_w73, 
            w74=> c0_n22_w74, 
            w75=> c0_n22_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n22_y
   );           
            
neuron_inst_23: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n23_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n23_w1, 
            w2=> c0_n23_w2, 
            w3=> c0_n23_w3, 
            w4=> c0_n23_w4, 
            w5=> c0_n23_w5, 
            w6=> c0_n23_w6, 
            w7=> c0_n23_w7, 
            w8=> c0_n23_w8, 
            w9=> c0_n23_w9, 
            w10=> c0_n23_w10, 
            w11=> c0_n23_w11, 
            w12=> c0_n23_w12, 
            w13=> c0_n23_w13, 
            w14=> c0_n23_w14, 
            w15=> c0_n23_w15, 
            w16=> c0_n23_w16, 
            w17=> c0_n23_w17, 
            w18=> c0_n23_w18, 
            w19=> c0_n23_w19, 
            w20=> c0_n23_w20, 
            w21=> c0_n23_w21, 
            w22=> c0_n23_w22, 
            w23=> c0_n23_w23, 
            w24=> c0_n23_w24, 
            w25=> c0_n23_w25, 
            w26=> c0_n23_w26, 
            w27=> c0_n23_w27, 
            w28=> c0_n23_w28, 
            w29=> c0_n23_w29, 
            w30=> c0_n23_w30, 
            w31=> c0_n23_w31, 
            w32=> c0_n23_w32, 
            w33=> c0_n23_w33, 
            w34=> c0_n23_w34, 
            w35=> c0_n23_w35, 
            w36=> c0_n23_w36, 
            w37=> c0_n23_w37, 
            w38=> c0_n23_w38, 
            w39=> c0_n23_w39, 
            w40=> c0_n23_w40, 
            w41=> c0_n23_w41, 
            w42=> c0_n23_w42, 
            w43=> c0_n23_w43, 
            w44=> c0_n23_w44, 
            w45=> c0_n23_w45, 
            w46=> c0_n23_w46, 
            w47=> c0_n23_w47, 
            w48=> c0_n23_w48, 
            w49=> c0_n23_w49, 
            w50=> c0_n23_w50, 
            w51=> c0_n23_w51, 
            w52=> c0_n23_w52, 
            w53=> c0_n23_w53, 
            w54=> c0_n23_w54, 
            w55=> c0_n23_w55, 
            w56=> c0_n23_w56, 
            w57=> c0_n23_w57, 
            w58=> c0_n23_w58, 
            w59=> c0_n23_w59, 
            w60=> c0_n23_w60, 
            w61=> c0_n23_w61, 
            w62=> c0_n23_w62, 
            w63=> c0_n23_w63, 
            w64=> c0_n23_w64, 
            w65=> c0_n23_w65, 
            w66=> c0_n23_w66, 
            w67=> c0_n23_w67, 
            w68=> c0_n23_w68, 
            w69=> c0_n23_w69, 
            w70=> c0_n23_w70, 
            w71=> c0_n23_w71, 
            w72=> c0_n23_w72, 
            w73=> c0_n23_w73, 
            w74=> c0_n23_w74, 
            w75=> c0_n23_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n23_y
   );           
            
neuron_inst_24: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n24_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n24_w1, 
            w2=> c0_n24_w2, 
            w3=> c0_n24_w3, 
            w4=> c0_n24_w4, 
            w5=> c0_n24_w5, 
            w6=> c0_n24_w6, 
            w7=> c0_n24_w7, 
            w8=> c0_n24_w8, 
            w9=> c0_n24_w9, 
            w10=> c0_n24_w10, 
            w11=> c0_n24_w11, 
            w12=> c0_n24_w12, 
            w13=> c0_n24_w13, 
            w14=> c0_n24_w14, 
            w15=> c0_n24_w15, 
            w16=> c0_n24_w16, 
            w17=> c0_n24_w17, 
            w18=> c0_n24_w18, 
            w19=> c0_n24_w19, 
            w20=> c0_n24_w20, 
            w21=> c0_n24_w21, 
            w22=> c0_n24_w22, 
            w23=> c0_n24_w23, 
            w24=> c0_n24_w24, 
            w25=> c0_n24_w25, 
            w26=> c0_n24_w26, 
            w27=> c0_n24_w27, 
            w28=> c0_n24_w28, 
            w29=> c0_n24_w29, 
            w30=> c0_n24_w30, 
            w31=> c0_n24_w31, 
            w32=> c0_n24_w32, 
            w33=> c0_n24_w33, 
            w34=> c0_n24_w34, 
            w35=> c0_n24_w35, 
            w36=> c0_n24_w36, 
            w37=> c0_n24_w37, 
            w38=> c0_n24_w38, 
            w39=> c0_n24_w39, 
            w40=> c0_n24_w40, 
            w41=> c0_n24_w41, 
            w42=> c0_n24_w42, 
            w43=> c0_n24_w43, 
            w44=> c0_n24_w44, 
            w45=> c0_n24_w45, 
            w46=> c0_n24_w46, 
            w47=> c0_n24_w47, 
            w48=> c0_n24_w48, 
            w49=> c0_n24_w49, 
            w50=> c0_n24_w50, 
            w51=> c0_n24_w51, 
            w52=> c0_n24_w52, 
            w53=> c0_n24_w53, 
            w54=> c0_n24_w54, 
            w55=> c0_n24_w55, 
            w56=> c0_n24_w56, 
            w57=> c0_n24_w57, 
            w58=> c0_n24_w58, 
            w59=> c0_n24_w59, 
            w60=> c0_n24_w60, 
            w61=> c0_n24_w61, 
            w62=> c0_n24_w62, 
            w63=> c0_n24_w63, 
            w64=> c0_n24_w64, 
            w65=> c0_n24_w65, 
            w66=> c0_n24_w66, 
            w67=> c0_n24_w67, 
            w68=> c0_n24_w68, 
            w69=> c0_n24_w69, 
            w70=> c0_n24_w70, 
            w71=> c0_n24_w71, 
            w72=> c0_n24_w72, 
            w73=> c0_n24_w73, 
            w74=> c0_n24_w74, 
            w75=> c0_n24_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n24_y
   );           
            
neuron_inst_25: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n25_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n25_w1, 
            w2=> c0_n25_w2, 
            w3=> c0_n25_w3, 
            w4=> c0_n25_w4, 
            w5=> c0_n25_w5, 
            w6=> c0_n25_w6, 
            w7=> c0_n25_w7, 
            w8=> c0_n25_w8, 
            w9=> c0_n25_w9, 
            w10=> c0_n25_w10, 
            w11=> c0_n25_w11, 
            w12=> c0_n25_w12, 
            w13=> c0_n25_w13, 
            w14=> c0_n25_w14, 
            w15=> c0_n25_w15, 
            w16=> c0_n25_w16, 
            w17=> c0_n25_w17, 
            w18=> c0_n25_w18, 
            w19=> c0_n25_w19, 
            w20=> c0_n25_w20, 
            w21=> c0_n25_w21, 
            w22=> c0_n25_w22, 
            w23=> c0_n25_w23, 
            w24=> c0_n25_w24, 
            w25=> c0_n25_w25, 
            w26=> c0_n25_w26, 
            w27=> c0_n25_w27, 
            w28=> c0_n25_w28, 
            w29=> c0_n25_w29, 
            w30=> c0_n25_w30, 
            w31=> c0_n25_w31, 
            w32=> c0_n25_w32, 
            w33=> c0_n25_w33, 
            w34=> c0_n25_w34, 
            w35=> c0_n25_w35, 
            w36=> c0_n25_w36, 
            w37=> c0_n25_w37, 
            w38=> c0_n25_w38, 
            w39=> c0_n25_w39, 
            w40=> c0_n25_w40, 
            w41=> c0_n25_w41, 
            w42=> c0_n25_w42, 
            w43=> c0_n25_w43, 
            w44=> c0_n25_w44, 
            w45=> c0_n25_w45, 
            w46=> c0_n25_w46, 
            w47=> c0_n25_w47, 
            w48=> c0_n25_w48, 
            w49=> c0_n25_w49, 
            w50=> c0_n25_w50, 
            w51=> c0_n25_w51, 
            w52=> c0_n25_w52, 
            w53=> c0_n25_w53, 
            w54=> c0_n25_w54, 
            w55=> c0_n25_w55, 
            w56=> c0_n25_w56, 
            w57=> c0_n25_w57, 
            w58=> c0_n25_w58, 
            w59=> c0_n25_w59, 
            w60=> c0_n25_w60, 
            w61=> c0_n25_w61, 
            w62=> c0_n25_w62, 
            w63=> c0_n25_w63, 
            w64=> c0_n25_w64, 
            w65=> c0_n25_w65, 
            w66=> c0_n25_w66, 
            w67=> c0_n25_w67, 
            w68=> c0_n25_w68, 
            w69=> c0_n25_w69, 
            w70=> c0_n25_w70, 
            w71=> c0_n25_w71, 
            w72=> c0_n25_w72, 
            w73=> c0_n25_w73, 
            w74=> c0_n25_w74, 
            w75=> c0_n25_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n25_y
   );           
            
neuron_inst_26: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n26_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n26_w1, 
            w2=> c0_n26_w2, 
            w3=> c0_n26_w3, 
            w4=> c0_n26_w4, 
            w5=> c0_n26_w5, 
            w6=> c0_n26_w6, 
            w7=> c0_n26_w7, 
            w8=> c0_n26_w8, 
            w9=> c0_n26_w9, 
            w10=> c0_n26_w10, 
            w11=> c0_n26_w11, 
            w12=> c0_n26_w12, 
            w13=> c0_n26_w13, 
            w14=> c0_n26_w14, 
            w15=> c0_n26_w15, 
            w16=> c0_n26_w16, 
            w17=> c0_n26_w17, 
            w18=> c0_n26_w18, 
            w19=> c0_n26_w19, 
            w20=> c0_n26_w20, 
            w21=> c0_n26_w21, 
            w22=> c0_n26_w22, 
            w23=> c0_n26_w23, 
            w24=> c0_n26_w24, 
            w25=> c0_n26_w25, 
            w26=> c0_n26_w26, 
            w27=> c0_n26_w27, 
            w28=> c0_n26_w28, 
            w29=> c0_n26_w29, 
            w30=> c0_n26_w30, 
            w31=> c0_n26_w31, 
            w32=> c0_n26_w32, 
            w33=> c0_n26_w33, 
            w34=> c0_n26_w34, 
            w35=> c0_n26_w35, 
            w36=> c0_n26_w36, 
            w37=> c0_n26_w37, 
            w38=> c0_n26_w38, 
            w39=> c0_n26_w39, 
            w40=> c0_n26_w40, 
            w41=> c0_n26_w41, 
            w42=> c0_n26_w42, 
            w43=> c0_n26_w43, 
            w44=> c0_n26_w44, 
            w45=> c0_n26_w45, 
            w46=> c0_n26_w46, 
            w47=> c0_n26_w47, 
            w48=> c0_n26_w48, 
            w49=> c0_n26_w49, 
            w50=> c0_n26_w50, 
            w51=> c0_n26_w51, 
            w52=> c0_n26_w52, 
            w53=> c0_n26_w53, 
            w54=> c0_n26_w54, 
            w55=> c0_n26_w55, 
            w56=> c0_n26_w56, 
            w57=> c0_n26_w57, 
            w58=> c0_n26_w58, 
            w59=> c0_n26_w59, 
            w60=> c0_n26_w60, 
            w61=> c0_n26_w61, 
            w62=> c0_n26_w62, 
            w63=> c0_n26_w63, 
            w64=> c0_n26_w64, 
            w65=> c0_n26_w65, 
            w66=> c0_n26_w66, 
            w67=> c0_n26_w67, 
            w68=> c0_n26_w68, 
            w69=> c0_n26_w69, 
            w70=> c0_n26_w70, 
            w71=> c0_n26_w71, 
            w72=> c0_n26_w72, 
            w73=> c0_n26_w73, 
            w74=> c0_n26_w74, 
            w75=> c0_n26_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n26_y
   );           
            
neuron_inst_27: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n27_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n27_w1, 
            w2=> c0_n27_w2, 
            w3=> c0_n27_w3, 
            w4=> c0_n27_w4, 
            w5=> c0_n27_w5, 
            w6=> c0_n27_w6, 
            w7=> c0_n27_w7, 
            w8=> c0_n27_w8, 
            w9=> c0_n27_w9, 
            w10=> c0_n27_w10, 
            w11=> c0_n27_w11, 
            w12=> c0_n27_w12, 
            w13=> c0_n27_w13, 
            w14=> c0_n27_w14, 
            w15=> c0_n27_w15, 
            w16=> c0_n27_w16, 
            w17=> c0_n27_w17, 
            w18=> c0_n27_w18, 
            w19=> c0_n27_w19, 
            w20=> c0_n27_w20, 
            w21=> c0_n27_w21, 
            w22=> c0_n27_w22, 
            w23=> c0_n27_w23, 
            w24=> c0_n27_w24, 
            w25=> c0_n27_w25, 
            w26=> c0_n27_w26, 
            w27=> c0_n27_w27, 
            w28=> c0_n27_w28, 
            w29=> c0_n27_w29, 
            w30=> c0_n27_w30, 
            w31=> c0_n27_w31, 
            w32=> c0_n27_w32, 
            w33=> c0_n27_w33, 
            w34=> c0_n27_w34, 
            w35=> c0_n27_w35, 
            w36=> c0_n27_w36, 
            w37=> c0_n27_w37, 
            w38=> c0_n27_w38, 
            w39=> c0_n27_w39, 
            w40=> c0_n27_w40, 
            w41=> c0_n27_w41, 
            w42=> c0_n27_w42, 
            w43=> c0_n27_w43, 
            w44=> c0_n27_w44, 
            w45=> c0_n27_w45, 
            w46=> c0_n27_w46, 
            w47=> c0_n27_w47, 
            w48=> c0_n27_w48, 
            w49=> c0_n27_w49, 
            w50=> c0_n27_w50, 
            w51=> c0_n27_w51, 
            w52=> c0_n27_w52, 
            w53=> c0_n27_w53, 
            w54=> c0_n27_w54, 
            w55=> c0_n27_w55, 
            w56=> c0_n27_w56, 
            w57=> c0_n27_w57, 
            w58=> c0_n27_w58, 
            w59=> c0_n27_w59, 
            w60=> c0_n27_w60, 
            w61=> c0_n27_w61, 
            w62=> c0_n27_w62, 
            w63=> c0_n27_w63, 
            w64=> c0_n27_w64, 
            w65=> c0_n27_w65, 
            w66=> c0_n27_w66, 
            w67=> c0_n27_w67, 
            w68=> c0_n27_w68, 
            w69=> c0_n27_w69, 
            w70=> c0_n27_w70, 
            w71=> c0_n27_w71, 
            w72=> c0_n27_w72, 
            w73=> c0_n27_w73, 
            w74=> c0_n27_w74, 
            w75=> c0_n27_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n27_y
   );           
            
neuron_inst_28: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n28_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n28_w1, 
            w2=> c0_n28_w2, 
            w3=> c0_n28_w3, 
            w4=> c0_n28_w4, 
            w5=> c0_n28_w5, 
            w6=> c0_n28_w6, 
            w7=> c0_n28_w7, 
            w8=> c0_n28_w8, 
            w9=> c0_n28_w9, 
            w10=> c0_n28_w10, 
            w11=> c0_n28_w11, 
            w12=> c0_n28_w12, 
            w13=> c0_n28_w13, 
            w14=> c0_n28_w14, 
            w15=> c0_n28_w15, 
            w16=> c0_n28_w16, 
            w17=> c0_n28_w17, 
            w18=> c0_n28_w18, 
            w19=> c0_n28_w19, 
            w20=> c0_n28_w20, 
            w21=> c0_n28_w21, 
            w22=> c0_n28_w22, 
            w23=> c0_n28_w23, 
            w24=> c0_n28_w24, 
            w25=> c0_n28_w25, 
            w26=> c0_n28_w26, 
            w27=> c0_n28_w27, 
            w28=> c0_n28_w28, 
            w29=> c0_n28_w29, 
            w30=> c0_n28_w30, 
            w31=> c0_n28_w31, 
            w32=> c0_n28_w32, 
            w33=> c0_n28_w33, 
            w34=> c0_n28_w34, 
            w35=> c0_n28_w35, 
            w36=> c0_n28_w36, 
            w37=> c0_n28_w37, 
            w38=> c0_n28_w38, 
            w39=> c0_n28_w39, 
            w40=> c0_n28_w40, 
            w41=> c0_n28_w41, 
            w42=> c0_n28_w42, 
            w43=> c0_n28_w43, 
            w44=> c0_n28_w44, 
            w45=> c0_n28_w45, 
            w46=> c0_n28_w46, 
            w47=> c0_n28_w47, 
            w48=> c0_n28_w48, 
            w49=> c0_n28_w49, 
            w50=> c0_n28_w50, 
            w51=> c0_n28_w51, 
            w52=> c0_n28_w52, 
            w53=> c0_n28_w53, 
            w54=> c0_n28_w54, 
            w55=> c0_n28_w55, 
            w56=> c0_n28_w56, 
            w57=> c0_n28_w57, 
            w58=> c0_n28_w58, 
            w59=> c0_n28_w59, 
            w60=> c0_n28_w60, 
            w61=> c0_n28_w61, 
            w62=> c0_n28_w62, 
            w63=> c0_n28_w63, 
            w64=> c0_n28_w64, 
            w65=> c0_n28_w65, 
            w66=> c0_n28_w66, 
            w67=> c0_n28_w67, 
            w68=> c0_n28_w68, 
            w69=> c0_n28_w69, 
            w70=> c0_n28_w70, 
            w71=> c0_n28_w71, 
            w72=> c0_n28_w72, 
            w73=> c0_n28_w73, 
            w74=> c0_n28_w74, 
            w75=> c0_n28_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n28_y
   );           
            
neuron_inst_29: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n29_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n29_w1, 
            w2=> c0_n29_w2, 
            w3=> c0_n29_w3, 
            w4=> c0_n29_w4, 
            w5=> c0_n29_w5, 
            w6=> c0_n29_w6, 
            w7=> c0_n29_w7, 
            w8=> c0_n29_w8, 
            w9=> c0_n29_w9, 
            w10=> c0_n29_w10, 
            w11=> c0_n29_w11, 
            w12=> c0_n29_w12, 
            w13=> c0_n29_w13, 
            w14=> c0_n29_w14, 
            w15=> c0_n29_w15, 
            w16=> c0_n29_w16, 
            w17=> c0_n29_w17, 
            w18=> c0_n29_w18, 
            w19=> c0_n29_w19, 
            w20=> c0_n29_w20, 
            w21=> c0_n29_w21, 
            w22=> c0_n29_w22, 
            w23=> c0_n29_w23, 
            w24=> c0_n29_w24, 
            w25=> c0_n29_w25, 
            w26=> c0_n29_w26, 
            w27=> c0_n29_w27, 
            w28=> c0_n29_w28, 
            w29=> c0_n29_w29, 
            w30=> c0_n29_w30, 
            w31=> c0_n29_w31, 
            w32=> c0_n29_w32, 
            w33=> c0_n29_w33, 
            w34=> c0_n29_w34, 
            w35=> c0_n29_w35, 
            w36=> c0_n29_w36, 
            w37=> c0_n29_w37, 
            w38=> c0_n29_w38, 
            w39=> c0_n29_w39, 
            w40=> c0_n29_w40, 
            w41=> c0_n29_w41, 
            w42=> c0_n29_w42, 
            w43=> c0_n29_w43, 
            w44=> c0_n29_w44, 
            w45=> c0_n29_w45, 
            w46=> c0_n29_w46, 
            w47=> c0_n29_w47, 
            w48=> c0_n29_w48, 
            w49=> c0_n29_w49, 
            w50=> c0_n29_w50, 
            w51=> c0_n29_w51, 
            w52=> c0_n29_w52, 
            w53=> c0_n29_w53, 
            w54=> c0_n29_w54, 
            w55=> c0_n29_w55, 
            w56=> c0_n29_w56, 
            w57=> c0_n29_w57, 
            w58=> c0_n29_w58, 
            w59=> c0_n29_w59, 
            w60=> c0_n29_w60, 
            w61=> c0_n29_w61, 
            w62=> c0_n29_w62, 
            w63=> c0_n29_w63, 
            w64=> c0_n29_w64, 
            w65=> c0_n29_w65, 
            w66=> c0_n29_w66, 
            w67=> c0_n29_w67, 
            w68=> c0_n29_w68, 
            w69=> c0_n29_w69, 
            w70=> c0_n29_w70, 
            w71=> c0_n29_w71, 
            w72=> c0_n29_w72, 
            w73=> c0_n29_w73, 
            w74=> c0_n29_w74, 
            w75=> c0_n29_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n29_y
   );           
            
neuron_inst_30: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n30_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n30_w1, 
            w2=> c0_n30_w2, 
            w3=> c0_n30_w3, 
            w4=> c0_n30_w4, 
            w5=> c0_n30_w5, 
            w6=> c0_n30_w6, 
            w7=> c0_n30_w7, 
            w8=> c0_n30_w8, 
            w9=> c0_n30_w9, 
            w10=> c0_n30_w10, 
            w11=> c0_n30_w11, 
            w12=> c0_n30_w12, 
            w13=> c0_n30_w13, 
            w14=> c0_n30_w14, 
            w15=> c0_n30_w15, 
            w16=> c0_n30_w16, 
            w17=> c0_n30_w17, 
            w18=> c0_n30_w18, 
            w19=> c0_n30_w19, 
            w20=> c0_n30_w20, 
            w21=> c0_n30_w21, 
            w22=> c0_n30_w22, 
            w23=> c0_n30_w23, 
            w24=> c0_n30_w24, 
            w25=> c0_n30_w25, 
            w26=> c0_n30_w26, 
            w27=> c0_n30_w27, 
            w28=> c0_n30_w28, 
            w29=> c0_n30_w29, 
            w30=> c0_n30_w30, 
            w31=> c0_n30_w31, 
            w32=> c0_n30_w32, 
            w33=> c0_n30_w33, 
            w34=> c0_n30_w34, 
            w35=> c0_n30_w35, 
            w36=> c0_n30_w36, 
            w37=> c0_n30_w37, 
            w38=> c0_n30_w38, 
            w39=> c0_n30_w39, 
            w40=> c0_n30_w40, 
            w41=> c0_n30_w41, 
            w42=> c0_n30_w42, 
            w43=> c0_n30_w43, 
            w44=> c0_n30_w44, 
            w45=> c0_n30_w45, 
            w46=> c0_n30_w46, 
            w47=> c0_n30_w47, 
            w48=> c0_n30_w48, 
            w49=> c0_n30_w49, 
            w50=> c0_n30_w50, 
            w51=> c0_n30_w51, 
            w52=> c0_n30_w52, 
            w53=> c0_n30_w53, 
            w54=> c0_n30_w54, 
            w55=> c0_n30_w55, 
            w56=> c0_n30_w56, 
            w57=> c0_n30_w57, 
            w58=> c0_n30_w58, 
            w59=> c0_n30_w59, 
            w60=> c0_n30_w60, 
            w61=> c0_n30_w61, 
            w62=> c0_n30_w62, 
            w63=> c0_n30_w63, 
            w64=> c0_n30_w64, 
            w65=> c0_n30_w65, 
            w66=> c0_n30_w66, 
            w67=> c0_n30_w67, 
            w68=> c0_n30_w68, 
            w69=> c0_n30_w69, 
            w70=> c0_n30_w70, 
            w71=> c0_n30_w71, 
            w72=> c0_n30_w72, 
            w73=> c0_n30_w73, 
            w74=> c0_n30_w74, 
            w75=> c0_n30_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n30_y
   );           
            
neuron_inst_31: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n31_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n31_w1, 
            w2=> c0_n31_w2, 
            w3=> c0_n31_w3, 
            w4=> c0_n31_w4, 
            w5=> c0_n31_w5, 
            w6=> c0_n31_w6, 
            w7=> c0_n31_w7, 
            w8=> c0_n31_w8, 
            w9=> c0_n31_w9, 
            w10=> c0_n31_w10, 
            w11=> c0_n31_w11, 
            w12=> c0_n31_w12, 
            w13=> c0_n31_w13, 
            w14=> c0_n31_w14, 
            w15=> c0_n31_w15, 
            w16=> c0_n31_w16, 
            w17=> c0_n31_w17, 
            w18=> c0_n31_w18, 
            w19=> c0_n31_w19, 
            w20=> c0_n31_w20, 
            w21=> c0_n31_w21, 
            w22=> c0_n31_w22, 
            w23=> c0_n31_w23, 
            w24=> c0_n31_w24, 
            w25=> c0_n31_w25, 
            w26=> c0_n31_w26, 
            w27=> c0_n31_w27, 
            w28=> c0_n31_w28, 
            w29=> c0_n31_w29, 
            w30=> c0_n31_w30, 
            w31=> c0_n31_w31, 
            w32=> c0_n31_w32, 
            w33=> c0_n31_w33, 
            w34=> c0_n31_w34, 
            w35=> c0_n31_w35, 
            w36=> c0_n31_w36, 
            w37=> c0_n31_w37, 
            w38=> c0_n31_w38, 
            w39=> c0_n31_w39, 
            w40=> c0_n31_w40, 
            w41=> c0_n31_w41, 
            w42=> c0_n31_w42, 
            w43=> c0_n31_w43, 
            w44=> c0_n31_w44, 
            w45=> c0_n31_w45, 
            w46=> c0_n31_w46, 
            w47=> c0_n31_w47, 
            w48=> c0_n31_w48, 
            w49=> c0_n31_w49, 
            w50=> c0_n31_w50, 
            w51=> c0_n31_w51, 
            w52=> c0_n31_w52, 
            w53=> c0_n31_w53, 
            w54=> c0_n31_w54, 
            w55=> c0_n31_w55, 
            w56=> c0_n31_w56, 
            w57=> c0_n31_w57, 
            w58=> c0_n31_w58, 
            w59=> c0_n31_w59, 
            w60=> c0_n31_w60, 
            w61=> c0_n31_w61, 
            w62=> c0_n31_w62, 
            w63=> c0_n31_w63, 
            w64=> c0_n31_w64, 
            w65=> c0_n31_w65, 
            w66=> c0_n31_w66, 
            w67=> c0_n31_w67, 
            w68=> c0_n31_w68, 
            w69=> c0_n31_w69, 
            w70=> c0_n31_w70, 
            w71=> c0_n31_w71, 
            w72=> c0_n31_w72, 
            w73=> c0_n31_w73, 
            w74=> c0_n31_w74, 
            w75=> c0_n31_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n31_y
   );           
            
neuron_inst_32: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n32_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n32_w1, 
            w2=> c0_n32_w2, 
            w3=> c0_n32_w3, 
            w4=> c0_n32_w4, 
            w5=> c0_n32_w5, 
            w6=> c0_n32_w6, 
            w7=> c0_n32_w7, 
            w8=> c0_n32_w8, 
            w9=> c0_n32_w9, 
            w10=> c0_n32_w10, 
            w11=> c0_n32_w11, 
            w12=> c0_n32_w12, 
            w13=> c0_n32_w13, 
            w14=> c0_n32_w14, 
            w15=> c0_n32_w15, 
            w16=> c0_n32_w16, 
            w17=> c0_n32_w17, 
            w18=> c0_n32_w18, 
            w19=> c0_n32_w19, 
            w20=> c0_n32_w20, 
            w21=> c0_n32_w21, 
            w22=> c0_n32_w22, 
            w23=> c0_n32_w23, 
            w24=> c0_n32_w24, 
            w25=> c0_n32_w25, 
            w26=> c0_n32_w26, 
            w27=> c0_n32_w27, 
            w28=> c0_n32_w28, 
            w29=> c0_n32_w29, 
            w30=> c0_n32_w30, 
            w31=> c0_n32_w31, 
            w32=> c0_n32_w32, 
            w33=> c0_n32_w33, 
            w34=> c0_n32_w34, 
            w35=> c0_n32_w35, 
            w36=> c0_n32_w36, 
            w37=> c0_n32_w37, 
            w38=> c0_n32_w38, 
            w39=> c0_n32_w39, 
            w40=> c0_n32_w40, 
            w41=> c0_n32_w41, 
            w42=> c0_n32_w42, 
            w43=> c0_n32_w43, 
            w44=> c0_n32_w44, 
            w45=> c0_n32_w45, 
            w46=> c0_n32_w46, 
            w47=> c0_n32_w47, 
            w48=> c0_n32_w48, 
            w49=> c0_n32_w49, 
            w50=> c0_n32_w50, 
            w51=> c0_n32_w51, 
            w52=> c0_n32_w52, 
            w53=> c0_n32_w53, 
            w54=> c0_n32_w54, 
            w55=> c0_n32_w55, 
            w56=> c0_n32_w56, 
            w57=> c0_n32_w57, 
            w58=> c0_n32_w58, 
            w59=> c0_n32_w59, 
            w60=> c0_n32_w60, 
            w61=> c0_n32_w61, 
            w62=> c0_n32_w62, 
            w63=> c0_n32_w63, 
            w64=> c0_n32_w64, 
            w65=> c0_n32_w65, 
            w66=> c0_n32_w66, 
            w67=> c0_n32_w67, 
            w68=> c0_n32_w68, 
            w69=> c0_n32_w69, 
            w70=> c0_n32_w70, 
            w71=> c0_n32_w71, 
            w72=> c0_n32_w72, 
            w73=> c0_n32_w73, 
            w74=> c0_n32_w74, 
            w75=> c0_n32_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n32_y
   );           
            
neuron_inst_33: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n33_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n33_w1, 
            w2=> c0_n33_w2, 
            w3=> c0_n33_w3, 
            w4=> c0_n33_w4, 
            w5=> c0_n33_w5, 
            w6=> c0_n33_w6, 
            w7=> c0_n33_w7, 
            w8=> c0_n33_w8, 
            w9=> c0_n33_w9, 
            w10=> c0_n33_w10, 
            w11=> c0_n33_w11, 
            w12=> c0_n33_w12, 
            w13=> c0_n33_w13, 
            w14=> c0_n33_w14, 
            w15=> c0_n33_w15, 
            w16=> c0_n33_w16, 
            w17=> c0_n33_w17, 
            w18=> c0_n33_w18, 
            w19=> c0_n33_w19, 
            w20=> c0_n33_w20, 
            w21=> c0_n33_w21, 
            w22=> c0_n33_w22, 
            w23=> c0_n33_w23, 
            w24=> c0_n33_w24, 
            w25=> c0_n33_w25, 
            w26=> c0_n33_w26, 
            w27=> c0_n33_w27, 
            w28=> c0_n33_w28, 
            w29=> c0_n33_w29, 
            w30=> c0_n33_w30, 
            w31=> c0_n33_w31, 
            w32=> c0_n33_w32, 
            w33=> c0_n33_w33, 
            w34=> c0_n33_w34, 
            w35=> c0_n33_w35, 
            w36=> c0_n33_w36, 
            w37=> c0_n33_w37, 
            w38=> c0_n33_w38, 
            w39=> c0_n33_w39, 
            w40=> c0_n33_w40, 
            w41=> c0_n33_w41, 
            w42=> c0_n33_w42, 
            w43=> c0_n33_w43, 
            w44=> c0_n33_w44, 
            w45=> c0_n33_w45, 
            w46=> c0_n33_w46, 
            w47=> c0_n33_w47, 
            w48=> c0_n33_w48, 
            w49=> c0_n33_w49, 
            w50=> c0_n33_w50, 
            w51=> c0_n33_w51, 
            w52=> c0_n33_w52, 
            w53=> c0_n33_w53, 
            w54=> c0_n33_w54, 
            w55=> c0_n33_w55, 
            w56=> c0_n33_w56, 
            w57=> c0_n33_w57, 
            w58=> c0_n33_w58, 
            w59=> c0_n33_w59, 
            w60=> c0_n33_w60, 
            w61=> c0_n33_w61, 
            w62=> c0_n33_w62, 
            w63=> c0_n33_w63, 
            w64=> c0_n33_w64, 
            w65=> c0_n33_w65, 
            w66=> c0_n33_w66, 
            w67=> c0_n33_w67, 
            w68=> c0_n33_w68, 
            w69=> c0_n33_w69, 
            w70=> c0_n33_w70, 
            w71=> c0_n33_w71, 
            w72=> c0_n33_w72, 
            w73=> c0_n33_w73, 
            w74=> c0_n33_w74, 
            w75=> c0_n33_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n33_y
   );           
            
neuron_inst_34: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n34_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n34_w1, 
            w2=> c0_n34_w2, 
            w3=> c0_n34_w3, 
            w4=> c0_n34_w4, 
            w5=> c0_n34_w5, 
            w6=> c0_n34_w6, 
            w7=> c0_n34_w7, 
            w8=> c0_n34_w8, 
            w9=> c0_n34_w9, 
            w10=> c0_n34_w10, 
            w11=> c0_n34_w11, 
            w12=> c0_n34_w12, 
            w13=> c0_n34_w13, 
            w14=> c0_n34_w14, 
            w15=> c0_n34_w15, 
            w16=> c0_n34_w16, 
            w17=> c0_n34_w17, 
            w18=> c0_n34_w18, 
            w19=> c0_n34_w19, 
            w20=> c0_n34_w20, 
            w21=> c0_n34_w21, 
            w22=> c0_n34_w22, 
            w23=> c0_n34_w23, 
            w24=> c0_n34_w24, 
            w25=> c0_n34_w25, 
            w26=> c0_n34_w26, 
            w27=> c0_n34_w27, 
            w28=> c0_n34_w28, 
            w29=> c0_n34_w29, 
            w30=> c0_n34_w30, 
            w31=> c0_n34_w31, 
            w32=> c0_n34_w32, 
            w33=> c0_n34_w33, 
            w34=> c0_n34_w34, 
            w35=> c0_n34_w35, 
            w36=> c0_n34_w36, 
            w37=> c0_n34_w37, 
            w38=> c0_n34_w38, 
            w39=> c0_n34_w39, 
            w40=> c0_n34_w40, 
            w41=> c0_n34_w41, 
            w42=> c0_n34_w42, 
            w43=> c0_n34_w43, 
            w44=> c0_n34_w44, 
            w45=> c0_n34_w45, 
            w46=> c0_n34_w46, 
            w47=> c0_n34_w47, 
            w48=> c0_n34_w48, 
            w49=> c0_n34_w49, 
            w50=> c0_n34_w50, 
            w51=> c0_n34_w51, 
            w52=> c0_n34_w52, 
            w53=> c0_n34_w53, 
            w54=> c0_n34_w54, 
            w55=> c0_n34_w55, 
            w56=> c0_n34_w56, 
            w57=> c0_n34_w57, 
            w58=> c0_n34_w58, 
            w59=> c0_n34_w59, 
            w60=> c0_n34_w60, 
            w61=> c0_n34_w61, 
            w62=> c0_n34_w62, 
            w63=> c0_n34_w63, 
            w64=> c0_n34_w64, 
            w65=> c0_n34_w65, 
            w66=> c0_n34_w66, 
            w67=> c0_n34_w67, 
            w68=> c0_n34_w68, 
            w69=> c0_n34_w69, 
            w70=> c0_n34_w70, 
            w71=> c0_n34_w71, 
            w72=> c0_n34_w72, 
            w73=> c0_n34_w73, 
            w74=> c0_n34_w74, 
            w75=> c0_n34_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n34_y
   );           
            
neuron_inst_35: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n35_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n35_w1, 
            w2=> c0_n35_w2, 
            w3=> c0_n35_w3, 
            w4=> c0_n35_w4, 
            w5=> c0_n35_w5, 
            w6=> c0_n35_w6, 
            w7=> c0_n35_w7, 
            w8=> c0_n35_w8, 
            w9=> c0_n35_w9, 
            w10=> c0_n35_w10, 
            w11=> c0_n35_w11, 
            w12=> c0_n35_w12, 
            w13=> c0_n35_w13, 
            w14=> c0_n35_w14, 
            w15=> c0_n35_w15, 
            w16=> c0_n35_w16, 
            w17=> c0_n35_w17, 
            w18=> c0_n35_w18, 
            w19=> c0_n35_w19, 
            w20=> c0_n35_w20, 
            w21=> c0_n35_w21, 
            w22=> c0_n35_w22, 
            w23=> c0_n35_w23, 
            w24=> c0_n35_w24, 
            w25=> c0_n35_w25, 
            w26=> c0_n35_w26, 
            w27=> c0_n35_w27, 
            w28=> c0_n35_w28, 
            w29=> c0_n35_w29, 
            w30=> c0_n35_w30, 
            w31=> c0_n35_w31, 
            w32=> c0_n35_w32, 
            w33=> c0_n35_w33, 
            w34=> c0_n35_w34, 
            w35=> c0_n35_w35, 
            w36=> c0_n35_w36, 
            w37=> c0_n35_w37, 
            w38=> c0_n35_w38, 
            w39=> c0_n35_w39, 
            w40=> c0_n35_w40, 
            w41=> c0_n35_w41, 
            w42=> c0_n35_w42, 
            w43=> c0_n35_w43, 
            w44=> c0_n35_w44, 
            w45=> c0_n35_w45, 
            w46=> c0_n35_w46, 
            w47=> c0_n35_w47, 
            w48=> c0_n35_w48, 
            w49=> c0_n35_w49, 
            w50=> c0_n35_w50, 
            w51=> c0_n35_w51, 
            w52=> c0_n35_w52, 
            w53=> c0_n35_w53, 
            w54=> c0_n35_w54, 
            w55=> c0_n35_w55, 
            w56=> c0_n35_w56, 
            w57=> c0_n35_w57, 
            w58=> c0_n35_w58, 
            w59=> c0_n35_w59, 
            w60=> c0_n35_w60, 
            w61=> c0_n35_w61, 
            w62=> c0_n35_w62, 
            w63=> c0_n35_w63, 
            w64=> c0_n35_w64, 
            w65=> c0_n35_w65, 
            w66=> c0_n35_w66, 
            w67=> c0_n35_w67, 
            w68=> c0_n35_w68, 
            w69=> c0_n35_w69, 
            w70=> c0_n35_w70, 
            w71=> c0_n35_w71, 
            w72=> c0_n35_w72, 
            w73=> c0_n35_w73, 
            w74=> c0_n35_w74, 
            w75=> c0_n35_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n35_y
   );           
            
neuron_inst_36: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n36_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n36_w1, 
            w2=> c0_n36_w2, 
            w3=> c0_n36_w3, 
            w4=> c0_n36_w4, 
            w5=> c0_n36_w5, 
            w6=> c0_n36_w6, 
            w7=> c0_n36_w7, 
            w8=> c0_n36_w8, 
            w9=> c0_n36_w9, 
            w10=> c0_n36_w10, 
            w11=> c0_n36_w11, 
            w12=> c0_n36_w12, 
            w13=> c0_n36_w13, 
            w14=> c0_n36_w14, 
            w15=> c0_n36_w15, 
            w16=> c0_n36_w16, 
            w17=> c0_n36_w17, 
            w18=> c0_n36_w18, 
            w19=> c0_n36_w19, 
            w20=> c0_n36_w20, 
            w21=> c0_n36_w21, 
            w22=> c0_n36_w22, 
            w23=> c0_n36_w23, 
            w24=> c0_n36_w24, 
            w25=> c0_n36_w25, 
            w26=> c0_n36_w26, 
            w27=> c0_n36_w27, 
            w28=> c0_n36_w28, 
            w29=> c0_n36_w29, 
            w30=> c0_n36_w30, 
            w31=> c0_n36_w31, 
            w32=> c0_n36_w32, 
            w33=> c0_n36_w33, 
            w34=> c0_n36_w34, 
            w35=> c0_n36_w35, 
            w36=> c0_n36_w36, 
            w37=> c0_n36_w37, 
            w38=> c0_n36_w38, 
            w39=> c0_n36_w39, 
            w40=> c0_n36_w40, 
            w41=> c0_n36_w41, 
            w42=> c0_n36_w42, 
            w43=> c0_n36_w43, 
            w44=> c0_n36_w44, 
            w45=> c0_n36_w45, 
            w46=> c0_n36_w46, 
            w47=> c0_n36_w47, 
            w48=> c0_n36_w48, 
            w49=> c0_n36_w49, 
            w50=> c0_n36_w50, 
            w51=> c0_n36_w51, 
            w52=> c0_n36_w52, 
            w53=> c0_n36_w53, 
            w54=> c0_n36_w54, 
            w55=> c0_n36_w55, 
            w56=> c0_n36_w56, 
            w57=> c0_n36_w57, 
            w58=> c0_n36_w58, 
            w59=> c0_n36_w59, 
            w60=> c0_n36_w60, 
            w61=> c0_n36_w61, 
            w62=> c0_n36_w62, 
            w63=> c0_n36_w63, 
            w64=> c0_n36_w64, 
            w65=> c0_n36_w65, 
            w66=> c0_n36_w66, 
            w67=> c0_n36_w67, 
            w68=> c0_n36_w68, 
            w69=> c0_n36_w69, 
            w70=> c0_n36_w70, 
            w71=> c0_n36_w71, 
            w72=> c0_n36_w72, 
            w73=> c0_n36_w73, 
            w74=> c0_n36_w74, 
            w75=> c0_n36_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n36_y
   );           
            
neuron_inst_37: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n37_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n37_w1, 
            w2=> c0_n37_w2, 
            w3=> c0_n37_w3, 
            w4=> c0_n37_w4, 
            w5=> c0_n37_w5, 
            w6=> c0_n37_w6, 
            w7=> c0_n37_w7, 
            w8=> c0_n37_w8, 
            w9=> c0_n37_w9, 
            w10=> c0_n37_w10, 
            w11=> c0_n37_w11, 
            w12=> c0_n37_w12, 
            w13=> c0_n37_w13, 
            w14=> c0_n37_w14, 
            w15=> c0_n37_w15, 
            w16=> c0_n37_w16, 
            w17=> c0_n37_w17, 
            w18=> c0_n37_w18, 
            w19=> c0_n37_w19, 
            w20=> c0_n37_w20, 
            w21=> c0_n37_w21, 
            w22=> c0_n37_w22, 
            w23=> c0_n37_w23, 
            w24=> c0_n37_w24, 
            w25=> c0_n37_w25, 
            w26=> c0_n37_w26, 
            w27=> c0_n37_w27, 
            w28=> c0_n37_w28, 
            w29=> c0_n37_w29, 
            w30=> c0_n37_w30, 
            w31=> c0_n37_w31, 
            w32=> c0_n37_w32, 
            w33=> c0_n37_w33, 
            w34=> c0_n37_w34, 
            w35=> c0_n37_w35, 
            w36=> c0_n37_w36, 
            w37=> c0_n37_w37, 
            w38=> c0_n37_w38, 
            w39=> c0_n37_w39, 
            w40=> c0_n37_w40, 
            w41=> c0_n37_w41, 
            w42=> c0_n37_w42, 
            w43=> c0_n37_w43, 
            w44=> c0_n37_w44, 
            w45=> c0_n37_w45, 
            w46=> c0_n37_w46, 
            w47=> c0_n37_w47, 
            w48=> c0_n37_w48, 
            w49=> c0_n37_w49, 
            w50=> c0_n37_w50, 
            w51=> c0_n37_w51, 
            w52=> c0_n37_w52, 
            w53=> c0_n37_w53, 
            w54=> c0_n37_w54, 
            w55=> c0_n37_w55, 
            w56=> c0_n37_w56, 
            w57=> c0_n37_w57, 
            w58=> c0_n37_w58, 
            w59=> c0_n37_w59, 
            w60=> c0_n37_w60, 
            w61=> c0_n37_w61, 
            w62=> c0_n37_w62, 
            w63=> c0_n37_w63, 
            w64=> c0_n37_w64, 
            w65=> c0_n37_w65, 
            w66=> c0_n37_w66, 
            w67=> c0_n37_w67, 
            w68=> c0_n37_w68, 
            w69=> c0_n37_w69, 
            w70=> c0_n37_w70, 
            w71=> c0_n37_w71, 
            w72=> c0_n37_w72, 
            w73=> c0_n37_w73, 
            w74=> c0_n37_w74, 
            w75=> c0_n37_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n37_y
   );           
            
neuron_inst_38: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n38_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n38_w1, 
            w2=> c0_n38_w2, 
            w3=> c0_n38_w3, 
            w4=> c0_n38_w4, 
            w5=> c0_n38_w5, 
            w6=> c0_n38_w6, 
            w7=> c0_n38_w7, 
            w8=> c0_n38_w8, 
            w9=> c0_n38_w9, 
            w10=> c0_n38_w10, 
            w11=> c0_n38_w11, 
            w12=> c0_n38_w12, 
            w13=> c0_n38_w13, 
            w14=> c0_n38_w14, 
            w15=> c0_n38_w15, 
            w16=> c0_n38_w16, 
            w17=> c0_n38_w17, 
            w18=> c0_n38_w18, 
            w19=> c0_n38_w19, 
            w20=> c0_n38_w20, 
            w21=> c0_n38_w21, 
            w22=> c0_n38_w22, 
            w23=> c0_n38_w23, 
            w24=> c0_n38_w24, 
            w25=> c0_n38_w25, 
            w26=> c0_n38_w26, 
            w27=> c0_n38_w27, 
            w28=> c0_n38_w28, 
            w29=> c0_n38_w29, 
            w30=> c0_n38_w30, 
            w31=> c0_n38_w31, 
            w32=> c0_n38_w32, 
            w33=> c0_n38_w33, 
            w34=> c0_n38_w34, 
            w35=> c0_n38_w35, 
            w36=> c0_n38_w36, 
            w37=> c0_n38_w37, 
            w38=> c0_n38_w38, 
            w39=> c0_n38_w39, 
            w40=> c0_n38_w40, 
            w41=> c0_n38_w41, 
            w42=> c0_n38_w42, 
            w43=> c0_n38_w43, 
            w44=> c0_n38_w44, 
            w45=> c0_n38_w45, 
            w46=> c0_n38_w46, 
            w47=> c0_n38_w47, 
            w48=> c0_n38_w48, 
            w49=> c0_n38_w49, 
            w50=> c0_n38_w50, 
            w51=> c0_n38_w51, 
            w52=> c0_n38_w52, 
            w53=> c0_n38_w53, 
            w54=> c0_n38_w54, 
            w55=> c0_n38_w55, 
            w56=> c0_n38_w56, 
            w57=> c0_n38_w57, 
            w58=> c0_n38_w58, 
            w59=> c0_n38_w59, 
            w60=> c0_n38_w60, 
            w61=> c0_n38_w61, 
            w62=> c0_n38_w62, 
            w63=> c0_n38_w63, 
            w64=> c0_n38_w64, 
            w65=> c0_n38_w65, 
            w66=> c0_n38_w66, 
            w67=> c0_n38_w67, 
            w68=> c0_n38_w68, 
            w69=> c0_n38_w69, 
            w70=> c0_n38_w70, 
            w71=> c0_n38_w71, 
            w72=> c0_n38_w72, 
            w73=> c0_n38_w73, 
            w74=> c0_n38_w74, 
            w75=> c0_n38_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n38_y
   );           
            
neuron_inst_39: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n39_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n39_w1, 
            w2=> c0_n39_w2, 
            w3=> c0_n39_w3, 
            w4=> c0_n39_w4, 
            w5=> c0_n39_w5, 
            w6=> c0_n39_w6, 
            w7=> c0_n39_w7, 
            w8=> c0_n39_w8, 
            w9=> c0_n39_w9, 
            w10=> c0_n39_w10, 
            w11=> c0_n39_w11, 
            w12=> c0_n39_w12, 
            w13=> c0_n39_w13, 
            w14=> c0_n39_w14, 
            w15=> c0_n39_w15, 
            w16=> c0_n39_w16, 
            w17=> c0_n39_w17, 
            w18=> c0_n39_w18, 
            w19=> c0_n39_w19, 
            w20=> c0_n39_w20, 
            w21=> c0_n39_w21, 
            w22=> c0_n39_w22, 
            w23=> c0_n39_w23, 
            w24=> c0_n39_w24, 
            w25=> c0_n39_w25, 
            w26=> c0_n39_w26, 
            w27=> c0_n39_w27, 
            w28=> c0_n39_w28, 
            w29=> c0_n39_w29, 
            w30=> c0_n39_w30, 
            w31=> c0_n39_w31, 
            w32=> c0_n39_w32, 
            w33=> c0_n39_w33, 
            w34=> c0_n39_w34, 
            w35=> c0_n39_w35, 
            w36=> c0_n39_w36, 
            w37=> c0_n39_w37, 
            w38=> c0_n39_w38, 
            w39=> c0_n39_w39, 
            w40=> c0_n39_w40, 
            w41=> c0_n39_w41, 
            w42=> c0_n39_w42, 
            w43=> c0_n39_w43, 
            w44=> c0_n39_w44, 
            w45=> c0_n39_w45, 
            w46=> c0_n39_w46, 
            w47=> c0_n39_w47, 
            w48=> c0_n39_w48, 
            w49=> c0_n39_w49, 
            w50=> c0_n39_w50, 
            w51=> c0_n39_w51, 
            w52=> c0_n39_w52, 
            w53=> c0_n39_w53, 
            w54=> c0_n39_w54, 
            w55=> c0_n39_w55, 
            w56=> c0_n39_w56, 
            w57=> c0_n39_w57, 
            w58=> c0_n39_w58, 
            w59=> c0_n39_w59, 
            w60=> c0_n39_w60, 
            w61=> c0_n39_w61, 
            w62=> c0_n39_w62, 
            w63=> c0_n39_w63, 
            w64=> c0_n39_w64, 
            w65=> c0_n39_w65, 
            w66=> c0_n39_w66, 
            w67=> c0_n39_w67, 
            w68=> c0_n39_w68, 
            w69=> c0_n39_w69, 
            w70=> c0_n39_w70, 
            w71=> c0_n39_w71, 
            w72=> c0_n39_w72, 
            w73=> c0_n39_w73, 
            w74=> c0_n39_w74, 
            w75=> c0_n39_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n39_y
   );           
            
neuron_inst_40: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n40_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n40_w1, 
            w2=> c0_n40_w2, 
            w3=> c0_n40_w3, 
            w4=> c0_n40_w4, 
            w5=> c0_n40_w5, 
            w6=> c0_n40_w6, 
            w7=> c0_n40_w7, 
            w8=> c0_n40_w8, 
            w9=> c0_n40_w9, 
            w10=> c0_n40_w10, 
            w11=> c0_n40_w11, 
            w12=> c0_n40_w12, 
            w13=> c0_n40_w13, 
            w14=> c0_n40_w14, 
            w15=> c0_n40_w15, 
            w16=> c0_n40_w16, 
            w17=> c0_n40_w17, 
            w18=> c0_n40_w18, 
            w19=> c0_n40_w19, 
            w20=> c0_n40_w20, 
            w21=> c0_n40_w21, 
            w22=> c0_n40_w22, 
            w23=> c0_n40_w23, 
            w24=> c0_n40_w24, 
            w25=> c0_n40_w25, 
            w26=> c0_n40_w26, 
            w27=> c0_n40_w27, 
            w28=> c0_n40_w28, 
            w29=> c0_n40_w29, 
            w30=> c0_n40_w30, 
            w31=> c0_n40_w31, 
            w32=> c0_n40_w32, 
            w33=> c0_n40_w33, 
            w34=> c0_n40_w34, 
            w35=> c0_n40_w35, 
            w36=> c0_n40_w36, 
            w37=> c0_n40_w37, 
            w38=> c0_n40_w38, 
            w39=> c0_n40_w39, 
            w40=> c0_n40_w40, 
            w41=> c0_n40_w41, 
            w42=> c0_n40_w42, 
            w43=> c0_n40_w43, 
            w44=> c0_n40_w44, 
            w45=> c0_n40_w45, 
            w46=> c0_n40_w46, 
            w47=> c0_n40_w47, 
            w48=> c0_n40_w48, 
            w49=> c0_n40_w49, 
            w50=> c0_n40_w50, 
            w51=> c0_n40_w51, 
            w52=> c0_n40_w52, 
            w53=> c0_n40_w53, 
            w54=> c0_n40_w54, 
            w55=> c0_n40_w55, 
            w56=> c0_n40_w56, 
            w57=> c0_n40_w57, 
            w58=> c0_n40_w58, 
            w59=> c0_n40_w59, 
            w60=> c0_n40_w60, 
            w61=> c0_n40_w61, 
            w62=> c0_n40_w62, 
            w63=> c0_n40_w63, 
            w64=> c0_n40_w64, 
            w65=> c0_n40_w65, 
            w66=> c0_n40_w66, 
            w67=> c0_n40_w67, 
            w68=> c0_n40_w68, 
            w69=> c0_n40_w69, 
            w70=> c0_n40_w70, 
            w71=> c0_n40_w71, 
            w72=> c0_n40_w72, 
            w73=> c0_n40_w73, 
            w74=> c0_n40_w74, 
            w75=> c0_n40_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n40_y
   );           
            
neuron_inst_41: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n41_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n41_w1, 
            w2=> c0_n41_w2, 
            w3=> c0_n41_w3, 
            w4=> c0_n41_w4, 
            w5=> c0_n41_w5, 
            w6=> c0_n41_w6, 
            w7=> c0_n41_w7, 
            w8=> c0_n41_w8, 
            w9=> c0_n41_w9, 
            w10=> c0_n41_w10, 
            w11=> c0_n41_w11, 
            w12=> c0_n41_w12, 
            w13=> c0_n41_w13, 
            w14=> c0_n41_w14, 
            w15=> c0_n41_w15, 
            w16=> c0_n41_w16, 
            w17=> c0_n41_w17, 
            w18=> c0_n41_w18, 
            w19=> c0_n41_w19, 
            w20=> c0_n41_w20, 
            w21=> c0_n41_w21, 
            w22=> c0_n41_w22, 
            w23=> c0_n41_w23, 
            w24=> c0_n41_w24, 
            w25=> c0_n41_w25, 
            w26=> c0_n41_w26, 
            w27=> c0_n41_w27, 
            w28=> c0_n41_w28, 
            w29=> c0_n41_w29, 
            w30=> c0_n41_w30, 
            w31=> c0_n41_w31, 
            w32=> c0_n41_w32, 
            w33=> c0_n41_w33, 
            w34=> c0_n41_w34, 
            w35=> c0_n41_w35, 
            w36=> c0_n41_w36, 
            w37=> c0_n41_w37, 
            w38=> c0_n41_w38, 
            w39=> c0_n41_w39, 
            w40=> c0_n41_w40, 
            w41=> c0_n41_w41, 
            w42=> c0_n41_w42, 
            w43=> c0_n41_w43, 
            w44=> c0_n41_w44, 
            w45=> c0_n41_w45, 
            w46=> c0_n41_w46, 
            w47=> c0_n41_w47, 
            w48=> c0_n41_w48, 
            w49=> c0_n41_w49, 
            w50=> c0_n41_w50, 
            w51=> c0_n41_w51, 
            w52=> c0_n41_w52, 
            w53=> c0_n41_w53, 
            w54=> c0_n41_w54, 
            w55=> c0_n41_w55, 
            w56=> c0_n41_w56, 
            w57=> c0_n41_w57, 
            w58=> c0_n41_w58, 
            w59=> c0_n41_w59, 
            w60=> c0_n41_w60, 
            w61=> c0_n41_w61, 
            w62=> c0_n41_w62, 
            w63=> c0_n41_w63, 
            w64=> c0_n41_w64, 
            w65=> c0_n41_w65, 
            w66=> c0_n41_w66, 
            w67=> c0_n41_w67, 
            w68=> c0_n41_w68, 
            w69=> c0_n41_w69, 
            w70=> c0_n41_w70, 
            w71=> c0_n41_w71, 
            w72=> c0_n41_w72, 
            w73=> c0_n41_w73, 
            w74=> c0_n41_w74, 
            w75=> c0_n41_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n41_y
   );           
            
neuron_inst_42: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n42_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n42_w1, 
            w2=> c0_n42_w2, 
            w3=> c0_n42_w3, 
            w4=> c0_n42_w4, 
            w5=> c0_n42_w5, 
            w6=> c0_n42_w6, 
            w7=> c0_n42_w7, 
            w8=> c0_n42_w8, 
            w9=> c0_n42_w9, 
            w10=> c0_n42_w10, 
            w11=> c0_n42_w11, 
            w12=> c0_n42_w12, 
            w13=> c0_n42_w13, 
            w14=> c0_n42_w14, 
            w15=> c0_n42_w15, 
            w16=> c0_n42_w16, 
            w17=> c0_n42_w17, 
            w18=> c0_n42_w18, 
            w19=> c0_n42_w19, 
            w20=> c0_n42_w20, 
            w21=> c0_n42_w21, 
            w22=> c0_n42_w22, 
            w23=> c0_n42_w23, 
            w24=> c0_n42_w24, 
            w25=> c0_n42_w25, 
            w26=> c0_n42_w26, 
            w27=> c0_n42_w27, 
            w28=> c0_n42_w28, 
            w29=> c0_n42_w29, 
            w30=> c0_n42_w30, 
            w31=> c0_n42_w31, 
            w32=> c0_n42_w32, 
            w33=> c0_n42_w33, 
            w34=> c0_n42_w34, 
            w35=> c0_n42_w35, 
            w36=> c0_n42_w36, 
            w37=> c0_n42_w37, 
            w38=> c0_n42_w38, 
            w39=> c0_n42_w39, 
            w40=> c0_n42_w40, 
            w41=> c0_n42_w41, 
            w42=> c0_n42_w42, 
            w43=> c0_n42_w43, 
            w44=> c0_n42_w44, 
            w45=> c0_n42_w45, 
            w46=> c0_n42_w46, 
            w47=> c0_n42_w47, 
            w48=> c0_n42_w48, 
            w49=> c0_n42_w49, 
            w50=> c0_n42_w50, 
            w51=> c0_n42_w51, 
            w52=> c0_n42_w52, 
            w53=> c0_n42_w53, 
            w54=> c0_n42_w54, 
            w55=> c0_n42_w55, 
            w56=> c0_n42_w56, 
            w57=> c0_n42_w57, 
            w58=> c0_n42_w58, 
            w59=> c0_n42_w59, 
            w60=> c0_n42_w60, 
            w61=> c0_n42_w61, 
            w62=> c0_n42_w62, 
            w63=> c0_n42_w63, 
            w64=> c0_n42_w64, 
            w65=> c0_n42_w65, 
            w66=> c0_n42_w66, 
            w67=> c0_n42_w67, 
            w68=> c0_n42_w68, 
            w69=> c0_n42_w69, 
            w70=> c0_n42_w70, 
            w71=> c0_n42_w71, 
            w72=> c0_n42_w72, 
            w73=> c0_n42_w73, 
            w74=> c0_n42_w74, 
            w75=> c0_n42_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n42_y
   );           
            
neuron_inst_43: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n43_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n43_w1, 
            w2=> c0_n43_w2, 
            w3=> c0_n43_w3, 
            w4=> c0_n43_w4, 
            w5=> c0_n43_w5, 
            w6=> c0_n43_w6, 
            w7=> c0_n43_w7, 
            w8=> c0_n43_w8, 
            w9=> c0_n43_w9, 
            w10=> c0_n43_w10, 
            w11=> c0_n43_w11, 
            w12=> c0_n43_w12, 
            w13=> c0_n43_w13, 
            w14=> c0_n43_w14, 
            w15=> c0_n43_w15, 
            w16=> c0_n43_w16, 
            w17=> c0_n43_w17, 
            w18=> c0_n43_w18, 
            w19=> c0_n43_w19, 
            w20=> c0_n43_w20, 
            w21=> c0_n43_w21, 
            w22=> c0_n43_w22, 
            w23=> c0_n43_w23, 
            w24=> c0_n43_w24, 
            w25=> c0_n43_w25, 
            w26=> c0_n43_w26, 
            w27=> c0_n43_w27, 
            w28=> c0_n43_w28, 
            w29=> c0_n43_w29, 
            w30=> c0_n43_w30, 
            w31=> c0_n43_w31, 
            w32=> c0_n43_w32, 
            w33=> c0_n43_w33, 
            w34=> c0_n43_w34, 
            w35=> c0_n43_w35, 
            w36=> c0_n43_w36, 
            w37=> c0_n43_w37, 
            w38=> c0_n43_w38, 
            w39=> c0_n43_w39, 
            w40=> c0_n43_w40, 
            w41=> c0_n43_w41, 
            w42=> c0_n43_w42, 
            w43=> c0_n43_w43, 
            w44=> c0_n43_w44, 
            w45=> c0_n43_w45, 
            w46=> c0_n43_w46, 
            w47=> c0_n43_w47, 
            w48=> c0_n43_w48, 
            w49=> c0_n43_w49, 
            w50=> c0_n43_w50, 
            w51=> c0_n43_w51, 
            w52=> c0_n43_w52, 
            w53=> c0_n43_w53, 
            w54=> c0_n43_w54, 
            w55=> c0_n43_w55, 
            w56=> c0_n43_w56, 
            w57=> c0_n43_w57, 
            w58=> c0_n43_w58, 
            w59=> c0_n43_w59, 
            w60=> c0_n43_w60, 
            w61=> c0_n43_w61, 
            w62=> c0_n43_w62, 
            w63=> c0_n43_w63, 
            w64=> c0_n43_w64, 
            w65=> c0_n43_w65, 
            w66=> c0_n43_w66, 
            w67=> c0_n43_w67, 
            w68=> c0_n43_w68, 
            w69=> c0_n43_w69, 
            w70=> c0_n43_w70, 
            w71=> c0_n43_w71, 
            w72=> c0_n43_w72, 
            w73=> c0_n43_w73, 
            w74=> c0_n43_w74, 
            w75=> c0_n43_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n43_y
   );           
            
neuron_inst_44: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n44_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n44_w1, 
            w2=> c0_n44_w2, 
            w3=> c0_n44_w3, 
            w4=> c0_n44_w4, 
            w5=> c0_n44_w5, 
            w6=> c0_n44_w6, 
            w7=> c0_n44_w7, 
            w8=> c0_n44_w8, 
            w9=> c0_n44_w9, 
            w10=> c0_n44_w10, 
            w11=> c0_n44_w11, 
            w12=> c0_n44_w12, 
            w13=> c0_n44_w13, 
            w14=> c0_n44_w14, 
            w15=> c0_n44_w15, 
            w16=> c0_n44_w16, 
            w17=> c0_n44_w17, 
            w18=> c0_n44_w18, 
            w19=> c0_n44_w19, 
            w20=> c0_n44_w20, 
            w21=> c0_n44_w21, 
            w22=> c0_n44_w22, 
            w23=> c0_n44_w23, 
            w24=> c0_n44_w24, 
            w25=> c0_n44_w25, 
            w26=> c0_n44_w26, 
            w27=> c0_n44_w27, 
            w28=> c0_n44_w28, 
            w29=> c0_n44_w29, 
            w30=> c0_n44_w30, 
            w31=> c0_n44_w31, 
            w32=> c0_n44_w32, 
            w33=> c0_n44_w33, 
            w34=> c0_n44_w34, 
            w35=> c0_n44_w35, 
            w36=> c0_n44_w36, 
            w37=> c0_n44_w37, 
            w38=> c0_n44_w38, 
            w39=> c0_n44_w39, 
            w40=> c0_n44_w40, 
            w41=> c0_n44_w41, 
            w42=> c0_n44_w42, 
            w43=> c0_n44_w43, 
            w44=> c0_n44_w44, 
            w45=> c0_n44_w45, 
            w46=> c0_n44_w46, 
            w47=> c0_n44_w47, 
            w48=> c0_n44_w48, 
            w49=> c0_n44_w49, 
            w50=> c0_n44_w50, 
            w51=> c0_n44_w51, 
            w52=> c0_n44_w52, 
            w53=> c0_n44_w53, 
            w54=> c0_n44_w54, 
            w55=> c0_n44_w55, 
            w56=> c0_n44_w56, 
            w57=> c0_n44_w57, 
            w58=> c0_n44_w58, 
            w59=> c0_n44_w59, 
            w60=> c0_n44_w60, 
            w61=> c0_n44_w61, 
            w62=> c0_n44_w62, 
            w63=> c0_n44_w63, 
            w64=> c0_n44_w64, 
            w65=> c0_n44_w65, 
            w66=> c0_n44_w66, 
            w67=> c0_n44_w67, 
            w68=> c0_n44_w68, 
            w69=> c0_n44_w69, 
            w70=> c0_n44_w70, 
            w71=> c0_n44_w71, 
            w72=> c0_n44_w72, 
            w73=> c0_n44_w73, 
            w74=> c0_n44_w74, 
            w75=> c0_n44_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n44_y
   );           
            
neuron_inst_45: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n45_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n45_w1, 
            w2=> c0_n45_w2, 
            w3=> c0_n45_w3, 
            w4=> c0_n45_w4, 
            w5=> c0_n45_w5, 
            w6=> c0_n45_w6, 
            w7=> c0_n45_w7, 
            w8=> c0_n45_w8, 
            w9=> c0_n45_w9, 
            w10=> c0_n45_w10, 
            w11=> c0_n45_w11, 
            w12=> c0_n45_w12, 
            w13=> c0_n45_w13, 
            w14=> c0_n45_w14, 
            w15=> c0_n45_w15, 
            w16=> c0_n45_w16, 
            w17=> c0_n45_w17, 
            w18=> c0_n45_w18, 
            w19=> c0_n45_w19, 
            w20=> c0_n45_w20, 
            w21=> c0_n45_w21, 
            w22=> c0_n45_w22, 
            w23=> c0_n45_w23, 
            w24=> c0_n45_w24, 
            w25=> c0_n45_w25, 
            w26=> c0_n45_w26, 
            w27=> c0_n45_w27, 
            w28=> c0_n45_w28, 
            w29=> c0_n45_w29, 
            w30=> c0_n45_w30, 
            w31=> c0_n45_w31, 
            w32=> c0_n45_w32, 
            w33=> c0_n45_w33, 
            w34=> c0_n45_w34, 
            w35=> c0_n45_w35, 
            w36=> c0_n45_w36, 
            w37=> c0_n45_w37, 
            w38=> c0_n45_w38, 
            w39=> c0_n45_w39, 
            w40=> c0_n45_w40, 
            w41=> c0_n45_w41, 
            w42=> c0_n45_w42, 
            w43=> c0_n45_w43, 
            w44=> c0_n45_w44, 
            w45=> c0_n45_w45, 
            w46=> c0_n45_w46, 
            w47=> c0_n45_w47, 
            w48=> c0_n45_w48, 
            w49=> c0_n45_w49, 
            w50=> c0_n45_w50, 
            w51=> c0_n45_w51, 
            w52=> c0_n45_w52, 
            w53=> c0_n45_w53, 
            w54=> c0_n45_w54, 
            w55=> c0_n45_w55, 
            w56=> c0_n45_w56, 
            w57=> c0_n45_w57, 
            w58=> c0_n45_w58, 
            w59=> c0_n45_w59, 
            w60=> c0_n45_w60, 
            w61=> c0_n45_w61, 
            w62=> c0_n45_w62, 
            w63=> c0_n45_w63, 
            w64=> c0_n45_w64, 
            w65=> c0_n45_w65, 
            w66=> c0_n45_w66, 
            w67=> c0_n45_w67, 
            w68=> c0_n45_w68, 
            w69=> c0_n45_w69, 
            w70=> c0_n45_w70, 
            w71=> c0_n45_w71, 
            w72=> c0_n45_w72, 
            w73=> c0_n45_w73, 
            w74=> c0_n45_w74, 
            w75=> c0_n45_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n45_y
   );           
            
neuron_inst_46: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n46_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n46_w1, 
            w2=> c0_n46_w2, 
            w3=> c0_n46_w3, 
            w4=> c0_n46_w4, 
            w5=> c0_n46_w5, 
            w6=> c0_n46_w6, 
            w7=> c0_n46_w7, 
            w8=> c0_n46_w8, 
            w9=> c0_n46_w9, 
            w10=> c0_n46_w10, 
            w11=> c0_n46_w11, 
            w12=> c0_n46_w12, 
            w13=> c0_n46_w13, 
            w14=> c0_n46_w14, 
            w15=> c0_n46_w15, 
            w16=> c0_n46_w16, 
            w17=> c0_n46_w17, 
            w18=> c0_n46_w18, 
            w19=> c0_n46_w19, 
            w20=> c0_n46_w20, 
            w21=> c0_n46_w21, 
            w22=> c0_n46_w22, 
            w23=> c0_n46_w23, 
            w24=> c0_n46_w24, 
            w25=> c0_n46_w25, 
            w26=> c0_n46_w26, 
            w27=> c0_n46_w27, 
            w28=> c0_n46_w28, 
            w29=> c0_n46_w29, 
            w30=> c0_n46_w30, 
            w31=> c0_n46_w31, 
            w32=> c0_n46_w32, 
            w33=> c0_n46_w33, 
            w34=> c0_n46_w34, 
            w35=> c0_n46_w35, 
            w36=> c0_n46_w36, 
            w37=> c0_n46_w37, 
            w38=> c0_n46_w38, 
            w39=> c0_n46_w39, 
            w40=> c0_n46_w40, 
            w41=> c0_n46_w41, 
            w42=> c0_n46_w42, 
            w43=> c0_n46_w43, 
            w44=> c0_n46_w44, 
            w45=> c0_n46_w45, 
            w46=> c0_n46_w46, 
            w47=> c0_n46_w47, 
            w48=> c0_n46_w48, 
            w49=> c0_n46_w49, 
            w50=> c0_n46_w50, 
            w51=> c0_n46_w51, 
            w52=> c0_n46_w52, 
            w53=> c0_n46_w53, 
            w54=> c0_n46_w54, 
            w55=> c0_n46_w55, 
            w56=> c0_n46_w56, 
            w57=> c0_n46_w57, 
            w58=> c0_n46_w58, 
            w59=> c0_n46_w59, 
            w60=> c0_n46_w60, 
            w61=> c0_n46_w61, 
            w62=> c0_n46_w62, 
            w63=> c0_n46_w63, 
            w64=> c0_n46_w64, 
            w65=> c0_n46_w65, 
            w66=> c0_n46_w66, 
            w67=> c0_n46_w67, 
            w68=> c0_n46_w68, 
            w69=> c0_n46_w69, 
            w70=> c0_n46_w70, 
            w71=> c0_n46_w71, 
            w72=> c0_n46_w72, 
            w73=> c0_n46_w73, 
            w74=> c0_n46_w74, 
            w75=> c0_n46_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n46_y
   );           
            
neuron_inst_47: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n47_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n47_w1, 
            w2=> c0_n47_w2, 
            w3=> c0_n47_w3, 
            w4=> c0_n47_w4, 
            w5=> c0_n47_w5, 
            w6=> c0_n47_w6, 
            w7=> c0_n47_w7, 
            w8=> c0_n47_w8, 
            w9=> c0_n47_w9, 
            w10=> c0_n47_w10, 
            w11=> c0_n47_w11, 
            w12=> c0_n47_w12, 
            w13=> c0_n47_w13, 
            w14=> c0_n47_w14, 
            w15=> c0_n47_w15, 
            w16=> c0_n47_w16, 
            w17=> c0_n47_w17, 
            w18=> c0_n47_w18, 
            w19=> c0_n47_w19, 
            w20=> c0_n47_w20, 
            w21=> c0_n47_w21, 
            w22=> c0_n47_w22, 
            w23=> c0_n47_w23, 
            w24=> c0_n47_w24, 
            w25=> c0_n47_w25, 
            w26=> c0_n47_w26, 
            w27=> c0_n47_w27, 
            w28=> c0_n47_w28, 
            w29=> c0_n47_w29, 
            w30=> c0_n47_w30, 
            w31=> c0_n47_w31, 
            w32=> c0_n47_w32, 
            w33=> c0_n47_w33, 
            w34=> c0_n47_w34, 
            w35=> c0_n47_w35, 
            w36=> c0_n47_w36, 
            w37=> c0_n47_w37, 
            w38=> c0_n47_w38, 
            w39=> c0_n47_w39, 
            w40=> c0_n47_w40, 
            w41=> c0_n47_w41, 
            w42=> c0_n47_w42, 
            w43=> c0_n47_w43, 
            w44=> c0_n47_w44, 
            w45=> c0_n47_w45, 
            w46=> c0_n47_w46, 
            w47=> c0_n47_w47, 
            w48=> c0_n47_w48, 
            w49=> c0_n47_w49, 
            w50=> c0_n47_w50, 
            w51=> c0_n47_w51, 
            w52=> c0_n47_w52, 
            w53=> c0_n47_w53, 
            w54=> c0_n47_w54, 
            w55=> c0_n47_w55, 
            w56=> c0_n47_w56, 
            w57=> c0_n47_w57, 
            w58=> c0_n47_w58, 
            w59=> c0_n47_w59, 
            w60=> c0_n47_w60, 
            w61=> c0_n47_w61, 
            w62=> c0_n47_w62, 
            w63=> c0_n47_w63, 
            w64=> c0_n47_w64, 
            w65=> c0_n47_w65, 
            w66=> c0_n47_w66, 
            w67=> c0_n47_w67, 
            w68=> c0_n47_w68, 
            w69=> c0_n47_w69, 
            w70=> c0_n47_w70, 
            w71=> c0_n47_w71, 
            w72=> c0_n47_w72, 
            w73=> c0_n47_w73, 
            w74=> c0_n47_w74, 
            w75=> c0_n47_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n47_y
   );           
            
neuron_inst_48: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n48_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n48_w1, 
            w2=> c0_n48_w2, 
            w3=> c0_n48_w3, 
            w4=> c0_n48_w4, 
            w5=> c0_n48_w5, 
            w6=> c0_n48_w6, 
            w7=> c0_n48_w7, 
            w8=> c0_n48_w8, 
            w9=> c0_n48_w9, 
            w10=> c0_n48_w10, 
            w11=> c0_n48_w11, 
            w12=> c0_n48_w12, 
            w13=> c0_n48_w13, 
            w14=> c0_n48_w14, 
            w15=> c0_n48_w15, 
            w16=> c0_n48_w16, 
            w17=> c0_n48_w17, 
            w18=> c0_n48_w18, 
            w19=> c0_n48_w19, 
            w20=> c0_n48_w20, 
            w21=> c0_n48_w21, 
            w22=> c0_n48_w22, 
            w23=> c0_n48_w23, 
            w24=> c0_n48_w24, 
            w25=> c0_n48_w25, 
            w26=> c0_n48_w26, 
            w27=> c0_n48_w27, 
            w28=> c0_n48_w28, 
            w29=> c0_n48_w29, 
            w30=> c0_n48_w30, 
            w31=> c0_n48_w31, 
            w32=> c0_n48_w32, 
            w33=> c0_n48_w33, 
            w34=> c0_n48_w34, 
            w35=> c0_n48_w35, 
            w36=> c0_n48_w36, 
            w37=> c0_n48_w37, 
            w38=> c0_n48_w38, 
            w39=> c0_n48_w39, 
            w40=> c0_n48_w40, 
            w41=> c0_n48_w41, 
            w42=> c0_n48_w42, 
            w43=> c0_n48_w43, 
            w44=> c0_n48_w44, 
            w45=> c0_n48_w45, 
            w46=> c0_n48_w46, 
            w47=> c0_n48_w47, 
            w48=> c0_n48_w48, 
            w49=> c0_n48_w49, 
            w50=> c0_n48_w50, 
            w51=> c0_n48_w51, 
            w52=> c0_n48_w52, 
            w53=> c0_n48_w53, 
            w54=> c0_n48_w54, 
            w55=> c0_n48_w55, 
            w56=> c0_n48_w56, 
            w57=> c0_n48_w57, 
            w58=> c0_n48_w58, 
            w59=> c0_n48_w59, 
            w60=> c0_n48_w60, 
            w61=> c0_n48_w61, 
            w62=> c0_n48_w62, 
            w63=> c0_n48_w63, 
            w64=> c0_n48_w64, 
            w65=> c0_n48_w65, 
            w66=> c0_n48_w66, 
            w67=> c0_n48_w67, 
            w68=> c0_n48_w68, 
            w69=> c0_n48_w69, 
            w70=> c0_n48_w70, 
            w71=> c0_n48_w71, 
            w72=> c0_n48_w72, 
            w73=> c0_n48_w73, 
            w74=> c0_n48_w74, 
            w75=> c0_n48_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n48_y
   );           
            
neuron_inst_49: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n49_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n49_w1, 
            w2=> c0_n49_w2, 
            w3=> c0_n49_w3, 
            w4=> c0_n49_w4, 
            w5=> c0_n49_w5, 
            w6=> c0_n49_w6, 
            w7=> c0_n49_w7, 
            w8=> c0_n49_w8, 
            w9=> c0_n49_w9, 
            w10=> c0_n49_w10, 
            w11=> c0_n49_w11, 
            w12=> c0_n49_w12, 
            w13=> c0_n49_w13, 
            w14=> c0_n49_w14, 
            w15=> c0_n49_w15, 
            w16=> c0_n49_w16, 
            w17=> c0_n49_w17, 
            w18=> c0_n49_w18, 
            w19=> c0_n49_w19, 
            w20=> c0_n49_w20, 
            w21=> c0_n49_w21, 
            w22=> c0_n49_w22, 
            w23=> c0_n49_w23, 
            w24=> c0_n49_w24, 
            w25=> c0_n49_w25, 
            w26=> c0_n49_w26, 
            w27=> c0_n49_w27, 
            w28=> c0_n49_w28, 
            w29=> c0_n49_w29, 
            w30=> c0_n49_w30, 
            w31=> c0_n49_w31, 
            w32=> c0_n49_w32, 
            w33=> c0_n49_w33, 
            w34=> c0_n49_w34, 
            w35=> c0_n49_w35, 
            w36=> c0_n49_w36, 
            w37=> c0_n49_w37, 
            w38=> c0_n49_w38, 
            w39=> c0_n49_w39, 
            w40=> c0_n49_w40, 
            w41=> c0_n49_w41, 
            w42=> c0_n49_w42, 
            w43=> c0_n49_w43, 
            w44=> c0_n49_w44, 
            w45=> c0_n49_w45, 
            w46=> c0_n49_w46, 
            w47=> c0_n49_w47, 
            w48=> c0_n49_w48, 
            w49=> c0_n49_w49, 
            w50=> c0_n49_w50, 
            w51=> c0_n49_w51, 
            w52=> c0_n49_w52, 
            w53=> c0_n49_w53, 
            w54=> c0_n49_w54, 
            w55=> c0_n49_w55, 
            w56=> c0_n49_w56, 
            w57=> c0_n49_w57, 
            w58=> c0_n49_w58, 
            w59=> c0_n49_w59, 
            w60=> c0_n49_w60, 
            w61=> c0_n49_w61, 
            w62=> c0_n49_w62, 
            w63=> c0_n49_w63, 
            w64=> c0_n49_w64, 
            w65=> c0_n49_w65, 
            w66=> c0_n49_w66, 
            w67=> c0_n49_w67, 
            w68=> c0_n49_w68, 
            w69=> c0_n49_w69, 
            w70=> c0_n49_w70, 
            w71=> c0_n49_w71, 
            w72=> c0_n49_w72, 
            w73=> c0_n49_w73, 
            w74=> c0_n49_w74, 
            w75=> c0_n49_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n49_y
   );           
            
neuron_inst_50: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n50_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n50_w1, 
            w2=> c0_n50_w2, 
            w3=> c0_n50_w3, 
            w4=> c0_n50_w4, 
            w5=> c0_n50_w5, 
            w6=> c0_n50_w6, 
            w7=> c0_n50_w7, 
            w8=> c0_n50_w8, 
            w9=> c0_n50_w9, 
            w10=> c0_n50_w10, 
            w11=> c0_n50_w11, 
            w12=> c0_n50_w12, 
            w13=> c0_n50_w13, 
            w14=> c0_n50_w14, 
            w15=> c0_n50_w15, 
            w16=> c0_n50_w16, 
            w17=> c0_n50_w17, 
            w18=> c0_n50_w18, 
            w19=> c0_n50_w19, 
            w20=> c0_n50_w20, 
            w21=> c0_n50_w21, 
            w22=> c0_n50_w22, 
            w23=> c0_n50_w23, 
            w24=> c0_n50_w24, 
            w25=> c0_n50_w25, 
            w26=> c0_n50_w26, 
            w27=> c0_n50_w27, 
            w28=> c0_n50_w28, 
            w29=> c0_n50_w29, 
            w30=> c0_n50_w30, 
            w31=> c0_n50_w31, 
            w32=> c0_n50_w32, 
            w33=> c0_n50_w33, 
            w34=> c0_n50_w34, 
            w35=> c0_n50_w35, 
            w36=> c0_n50_w36, 
            w37=> c0_n50_w37, 
            w38=> c0_n50_w38, 
            w39=> c0_n50_w39, 
            w40=> c0_n50_w40, 
            w41=> c0_n50_w41, 
            w42=> c0_n50_w42, 
            w43=> c0_n50_w43, 
            w44=> c0_n50_w44, 
            w45=> c0_n50_w45, 
            w46=> c0_n50_w46, 
            w47=> c0_n50_w47, 
            w48=> c0_n50_w48, 
            w49=> c0_n50_w49, 
            w50=> c0_n50_w50, 
            w51=> c0_n50_w51, 
            w52=> c0_n50_w52, 
            w53=> c0_n50_w53, 
            w54=> c0_n50_w54, 
            w55=> c0_n50_w55, 
            w56=> c0_n50_w56, 
            w57=> c0_n50_w57, 
            w58=> c0_n50_w58, 
            w59=> c0_n50_w59, 
            w60=> c0_n50_w60, 
            w61=> c0_n50_w61, 
            w62=> c0_n50_w62, 
            w63=> c0_n50_w63, 
            w64=> c0_n50_w64, 
            w65=> c0_n50_w65, 
            w66=> c0_n50_w66, 
            w67=> c0_n50_w67, 
            w68=> c0_n50_w68, 
            w69=> c0_n50_w69, 
            w70=> c0_n50_w70, 
            w71=> c0_n50_w71, 
            w72=> c0_n50_w72, 
            w73=> c0_n50_w73, 
            w74=> c0_n50_w74, 
            w75=> c0_n50_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n50_y
   );           
            
neuron_inst_51: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n51_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n51_w1, 
            w2=> c0_n51_w2, 
            w3=> c0_n51_w3, 
            w4=> c0_n51_w4, 
            w5=> c0_n51_w5, 
            w6=> c0_n51_w6, 
            w7=> c0_n51_w7, 
            w8=> c0_n51_w8, 
            w9=> c0_n51_w9, 
            w10=> c0_n51_w10, 
            w11=> c0_n51_w11, 
            w12=> c0_n51_w12, 
            w13=> c0_n51_w13, 
            w14=> c0_n51_w14, 
            w15=> c0_n51_w15, 
            w16=> c0_n51_w16, 
            w17=> c0_n51_w17, 
            w18=> c0_n51_w18, 
            w19=> c0_n51_w19, 
            w20=> c0_n51_w20, 
            w21=> c0_n51_w21, 
            w22=> c0_n51_w22, 
            w23=> c0_n51_w23, 
            w24=> c0_n51_w24, 
            w25=> c0_n51_w25, 
            w26=> c0_n51_w26, 
            w27=> c0_n51_w27, 
            w28=> c0_n51_w28, 
            w29=> c0_n51_w29, 
            w30=> c0_n51_w30, 
            w31=> c0_n51_w31, 
            w32=> c0_n51_w32, 
            w33=> c0_n51_w33, 
            w34=> c0_n51_w34, 
            w35=> c0_n51_w35, 
            w36=> c0_n51_w36, 
            w37=> c0_n51_w37, 
            w38=> c0_n51_w38, 
            w39=> c0_n51_w39, 
            w40=> c0_n51_w40, 
            w41=> c0_n51_w41, 
            w42=> c0_n51_w42, 
            w43=> c0_n51_w43, 
            w44=> c0_n51_w44, 
            w45=> c0_n51_w45, 
            w46=> c0_n51_w46, 
            w47=> c0_n51_w47, 
            w48=> c0_n51_w48, 
            w49=> c0_n51_w49, 
            w50=> c0_n51_w50, 
            w51=> c0_n51_w51, 
            w52=> c0_n51_w52, 
            w53=> c0_n51_w53, 
            w54=> c0_n51_w54, 
            w55=> c0_n51_w55, 
            w56=> c0_n51_w56, 
            w57=> c0_n51_w57, 
            w58=> c0_n51_w58, 
            w59=> c0_n51_w59, 
            w60=> c0_n51_w60, 
            w61=> c0_n51_w61, 
            w62=> c0_n51_w62, 
            w63=> c0_n51_w63, 
            w64=> c0_n51_w64, 
            w65=> c0_n51_w65, 
            w66=> c0_n51_w66, 
            w67=> c0_n51_w67, 
            w68=> c0_n51_w68, 
            w69=> c0_n51_w69, 
            w70=> c0_n51_w70, 
            w71=> c0_n51_w71, 
            w72=> c0_n51_w72, 
            w73=> c0_n51_w73, 
            w74=> c0_n51_w74, 
            w75=> c0_n51_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n51_y
   );           
            
neuron_inst_52: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n52_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n52_w1, 
            w2=> c0_n52_w2, 
            w3=> c0_n52_w3, 
            w4=> c0_n52_w4, 
            w5=> c0_n52_w5, 
            w6=> c0_n52_w6, 
            w7=> c0_n52_w7, 
            w8=> c0_n52_w8, 
            w9=> c0_n52_w9, 
            w10=> c0_n52_w10, 
            w11=> c0_n52_w11, 
            w12=> c0_n52_w12, 
            w13=> c0_n52_w13, 
            w14=> c0_n52_w14, 
            w15=> c0_n52_w15, 
            w16=> c0_n52_w16, 
            w17=> c0_n52_w17, 
            w18=> c0_n52_w18, 
            w19=> c0_n52_w19, 
            w20=> c0_n52_w20, 
            w21=> c0_n52_w21, 
            w22=> c0_n52_w22, 
            w23=> c0_n52_w23, 
            w24=> c0_n52_w24, 
            w25=> c0_n52_w25, 
            w26=> c0_n52_w26, 
            w27=> c0_n52_w27, 
            w28=> c0_n52_w28, 
            w29=> c0_n52_w29, 
            w30=> c0_n52_w30, 
            w31=> c0_n52_w31, 
            w32=> c0_n52_w32, 
            w33=> c0_n52_w33, 
            w34=> c0_n52_w34, 
            w35=> c0_n52_w35, 
            w36=> c0_n52_w36, 
            w37=> c0_n52_w37, 
            w38=> c0_n52_w38, 
            w39=> c0_n52_w39, 
            w40=> c0_n52_w40, 
            w41=> c0_n52_w41, 
            w42=> c0_n52_w42, 
            w43=> c0_n52_w43, 
            w44=> c0_n52_w44, 
            w45=> c0_n52_w45, 
            w46=> c0_n52_w46, 
            w47=> c0_n52_w47, 
            w48=> c0_n52_w48, 
            w49=> c0_n52_w49, 
            w50=> c0_n52_w50, 
            w51=> c0_n52_w51, 
            w52=> c0_n52_w52, 
            w53=> c0_n52_w53, 
            w54=> c0_n52_w54, 
            w55=> c0_n52_w55, 
            w56=> c0_n52_w56, 
            w57=> c0_n52_w57, 
            w58=> c0_n52_w58, 
            w59=> c0_n52_w59, 
            w60=> c0_n52_w60, 
            w61=> c0_n52_w61, 
            w62=> c0_n52_w62, 
            w63=> c0_n52_w63, 
            w64=> c0_n52_w64, 
            w65=> c0_n52_w65, 
            w66=> c0_n52_w66, 
            w67=> c0_n52_w67, 
            w68=> c0_n52_w68, 
            w69=> c0_n52_w69, 
            w70=> c0_n52_w70, 
            w71=> c0_n52_w71, 
            w72=> c0_n52_w72, 
            w73=> c0_n52_w73, 
            w74=> c0_n52_w74, 
            w75=> c0_n52_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n52_y
   );           
            
neuron_inst_53: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n53_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n53_w1, 
            w2=> c0_n53_w2, 
            w3=> c0_n53_w3, 
            w4=> c0_n53_w4, 
            w5=> c0_n53_w5, 
            w6=> c0_n53_w6, 
            w7=> c0_n53_w7, 
            w8=> c0_n53_w8, 
            w9=> c0_n53_w9, 
            w10=> c0_n53_w10, 
            w11=> c0_n53_w11, 
            w12=> c0_n53_w12, 
            w13=> c0_n53_w13, 
            w14=> c0_n53_w14, 
            w15=> c0_n53_w15, 
            w16=> c0_n53_w16, 
            w17=> c0_n53_w17, 
            w18=> c0_n53_w18, 
            w19=> c0_n53_w19, 
            w20=> c0_n53_w20, 
            w21=> c0_n53_w21, 
            w22=> c0_n53_w22, 
            w23=> c0_n53_w23, 
            w24=> c0_n53_w24, 
            w25=> c0_n53_w25, 
            w26=> c0_n53_w26, 
            w27=> c0_n53_w27, 
            w28=> c0_n53_w28, 
            w29=> c0_n53_w29, 
            w30=> c0_n53_w30, 
            w31=> c0_n53_w31, 
            w32=> c0_n53_w32, 
            w33=> c0_n53_w33, 
            w34=> c0_n53_w34, 
            w35=> c0_n53_w35, 
            w36=> c0_n53_w36, 
            w37=> c0_n53_w37, 
            w38=> c0_n53_w38, 
            w39=> c0_n53_w39, 
            w40=> c0_n53_w40, 
            w41=> c0_n53_w41, 
            w42=> c0_n53_w42, 
            w43=> c0_n53_w43, 
            w44=> c0_n53_w44, 
            w45=> c0_n53_w45, 
            w46=> c0_n53_w46, 
            w47=> c0_n53_w47, 
            w48=> c0_n53_w48, 
            w49=> c0_n53_w49, 
            w50=> c0_n53_w50, 
            w51=> c0_n53_w51, 
            w52=> c0_n53_w52, 
            w53=> c0_n53_w53, 
            w54=> c0_n53_w54, 
            w55=> c0_n53_w55, 
            w56=> c0_n53_w56, 
            w57=> c0_n53_w57, 
            w58=> c0_n53_w58, 
            w59=> c0_n53_w59, 
            w60=> c0_n53_w60, 
            w61=> c0_n53_w61, 
            w62=> c0_n53_w62, 
            w63=> c0_n53_w63, 
            w64=> c0_n53_w64, 
            w65=> c0_n53_w65, 
            w66=> c0_n53_w66, 
            w67=> c0_n53_w67, 
            w68=> c0_n53_w68, 
            w69=> c0_n53_w69, 
            w70=> c0_n53_w70, 
            w71=> c0_n53_w71, 
            w72=> c0_n53_w72, 
            w73=> c0_n53_w73, 
            w74=> c0_n53_w74, 
            w75=> c0_n53_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n53_y
   );           
            
neuron_inst_54: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n54_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n54_w1, 
            w2=> c0_n54_w2, 
            w3=> c0_n54_w3, 
            w4=> c0_n54_w4, 
            w5=> c0_n54_w5, 
            w6=> c0_n54_w6, 
            w7=> c0_n54_w7, 
            w8=> c0_n54_w8, 
            w9=> c0_n54_w9, 
            w10=> c0_n54_w10, 
            w11=> c0_n54_w11, 
            w12=> c0_n54_w12, 
            w13=> c0_n54_w13, 
            w14=> c0_n54_w14, 
            w15=> c0_n54_w15, 
            w16=> c0_n54_w16, 
            w17=> c0_n54_w17, 
            w18=> c0_n54_w18, 
            w19=> c0_n54_w19, 
            w20=> c0_n54_w20, 
            w21=> c0_n54_w21, 
            w22=> c0_n54_w22, 
            w23=> c0_n54_w23, 
            w24=> c0_n54_w24, 
            w25=> c0_n54_w25, 
            w26=> c0_n54_w26, 
            w27=> c0_n54_w27, 
            w28=> c0_n54_w28, 
            w29=> c0_n54_w29, 
            w30=> c0_n54_w30, 
            w31=> c0_n54_w31, 
            w32=> c0_n54_w32, 
            w33=> c0_n54_w33, 
            w34=> c0_n54_w34, 
            w35=> c0_n54_w35, 
            w36=> c0_n54_w36, 
            w37=> c0_n54_w37, 
            w38=> c0_n54_w38, 
            w39=> c0_n54_w39, 
            w40=> c0_n54_w40, 
            w41=> c0_n54_w41, 
            w42=> c0_n54_w42, 
            w43=> c0_n54_w43, 
            w44=> c0_n54_w44, 
            w45=> c0_n54_w45, 
            w46=> c0_n54_w46, 
            w47=> c0_n54_w47, 
            w48=> c0_n54_w48, 
            w49=> c0_n54_w49, 
            w50=> c0_n54_w50, 
            w51=> c0_n54_w51, 
            w52=> c0_n54_w52, 
            w53=> c0_n54_w53, 
            w54=> c0_n54_w54, 
            w55=> c0_n54_w55, 
            w56=> c0_n54_w56, 
            w57=> c0_n54_w57, 
            w58=> c0_n54_w58, 
            w59=> c0_n54_w59, 
            w60=> c0_n54_w60, 
            w61=> c0_n54_w61, 
            w62=> c0_n54_w62, 
            w63=> c0_n54_w63, 
            w64=> c0_n54_w64, 
            w65=> c0_n54_w65, 
            w66=> c0_n54_w66, 
            w67=> c0_n54_w67, 
            w68=> c0_n54_w68, 
            w69=> c0_n54_w69, 
            w70=> c0_n54_w70, 
            w71=> c0_n54_w71, 
            w72=> c0_n54_w72, 
            w73=> c0_n54_w73, 
            w74=> c0_n54_w74, 
            w75=> c0_n54_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n54_y
   );           
            
neuron_inst_55: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n55_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n55_w1, 
            w2=> c0_n55_w2, 
            w3=> c0_n55_w3, 
            w4=> c0_n55_w4, 
            w5=> c0_n55_w5, 
            w6=> c0_n55_w6, 
            w7=> c0_n55_w7, 
            w8=> c0_n55_w8, 
            w9=> c0_n55_w9, 
            w10=> c0_n55_w10, 
            w11=> c0_n55_w11, 
            w12=> c0_n55_w12, 
            w13=> c0_n55_w13, 
            w14=> c0_n55_w14, 
            w15=> c0_n55_w15, 
            w16=> c0_n55_w16, 
            w17=> c0_n55_w17, 
            w18=> c0_n55_w18, 
            w19=> c0_n55_w19, 
            w20=> c0_n55_w20, 
            w21=> c0_n55_w21, 
            w22=> c0_n55_w22, 
            w23=> c0_n55_w23, 
            w24=> c0_n55_w24, 
            w25=> c0_n55_w25, 
            w26=> c0_n55_w26, 
            w27=> c0_n55_w27, 
            w28=> c0_n55_w28, 
            w29=> c0_n55_w29, 
            w30=> c0_n55_w30, 
            w31=> c0_n55_w31, 
            w32=> c0_n55_w32, 
            w33=> c0_n55_w33, 
            w34=> c0_n55_w34, 
            w35=> c0_n55_w35, 
            w36=> c0_n55_w36, 
            w37=> c0_n55_w37, 
            w38=> c0_n55_w38, 
            w39=> c0_n55_w39, 
            w40=> c0_n55_w40, 
            w41=> c0_n55_w41, 
            w42=> c0_n55_w42, 
            w43=> c0_n55_w43, 
            w44=> c0_n55_w44, 
            w45=> c0_n55_w45, 
            w46=> c0_n55_w46, 
            w47=> c0_n55_w47, 
            w48=> c0_n55_w48, 
            w49=> c0_n55_w49, 
            w50=> c0_n55_w50, 
            w51=> c0_n55_w51, 
            w52=> c0_n55_w52, 
            w53=> c0_n55_w53, 
            w54=> c0_n55_w54, 
            w55=> c0_n55_w55, 
            w56=> c0_n55_w56, 
            w57=> c0_n55_w57, 
            w58=> c0_n55_w58, 
            w59=> c0_n55_w59, 
            w60=> c0_n55_w60, 
            w61=> c0_n55_w61, 
            w62=> c0_n55_w62, 
            w63=> c0_n55_w63, 
            w64=> c0_n55_w64, 
            w65=> c0_n55_w65, 
            w66=> c0_n55_w66, 
            w67=> c0_n55_w67, 
            w68=> c0_n55_w68, 
            w69=> c0_n55_w69, 
            w70=> c0_n55_w70, 
            w71=> c0_n55_w71, 
            w72=> c0_n55_w72, 
            w73=> c0_n55_w73, 
            w74=> c0_n55_w74, 
            w75=> c0_n55_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n55_y
   );           
            
neuron_inst_56: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n56_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n56_w1, 
            w2=> c0_n56_w2, 
            w3=> c0_n56_w3, 
            w4=> c0_n56_w4, 
            w5=> c0_n56_w5, 
            w6=> c0_n56_w6, 
            w7=> c0_n56_w7, 
            w8=> c0_n56_w8, 
            w9=> c0_n56_w9, 
            w10=> c0_n56_w10, 
            w11=> c0_n56_w11, 
            w12=> c0_n56_w12, 
            w13=> c0_n56_w13, 
            w14=> c0_n56_w14, 
            w15=> c0_n56_w15, 
            w16=> c0_n56_w16, 
            w17=> c0_n56_w17, 
            w18=> c0_n56_w18, 
            w19=> c0_n56_w19, 
            w20=> c0_n56_w20, 
            w21=> c0_n56_w21, 
            w22=> c0_n56_w22, 
            w23=> c0_n56_w23, 
            w24=> c0_n56_w24, 
            w25=> c0_n56_w25, 
            w26=> c0_n56_w26, 
            w27=> c0_n56_w27, 
            w28=> c0_n56_w28, 
            w29=> c0_n56_w29, 
            w30=> c0_n56_w30, 
            w31=> c0_n56_w31, 
            w32=> c0_n56_w32, 
            w33=> c0_n56_w33, 
            w34=> c0_n56_w34, 
            w35=> c0_n56_w35, 
            w36=> c0_n56_w36, 
            w37=> c0_n56_w37, 
            w38=> c0_n56_w38, 
            w39=> c0_n56_w39, 
            w40=> c0_n56_w40, 
            w41=> c0_n56_w41, 
            w42=> c0_n56_w42, 
            w43=> c0_n56_w43, 
            w44=> c0_n56_w44, 
            w45=> c0_n56_w45, 
            w46=> c0_n56_w46, 
            w47=> c0_n56_w47, 
            w48=> c0_n56_w48, 
            w49=> c0_n56_w49, 
            w50=> c0_n56_w50, 
            w51=> c0_n56_w51, 
            w52=> c0_n56_w52, 
            w53=> c0_n56_w53, 
            w54=> c0_n56_w54, 
            w55=> c0_n56_w55, 
            w56=> c0_n56_w56, 
            w57=> c0_n56_w57, 
            w58=> c0_n56_w58, 
            w59=> c0_n56_w59, 
            w60=> c0_n56_w60, 
            w61=> c0_n56_w61, 
            w62=> c0_n56_w62, 
            w63=> c0_n56_w63, 
            w64=> c0_n56_w64, 
            w65=> c0_n56_w65, 
            w66=> c0_n56_w66, 
            w67=> c0_n56_w67, 
            w68=> c0_n56_w68, 
            w69=> c0_n56_w69, 
            w70=> c0_n56_w70, 
            w71=> c0_n56_w71, 
            w72=> c0_n56_w72, 
            w73=> c0_n56_w73, 
            w74=> c0_n56_w74, 
            w75=> c0_n56_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n56_y
   );           
            
neuron_inst_57: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n57_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n57_w1, 
            w2=> c0_n57_w2, 
            w3=> c0_n57_w3, 
            w4=> c0_n57_w4, 
            w5=> c0_n57_w5, 
            w6=> c0_n57_w6, 
            w7=> c0_n57_w7, 
            w8=> c0_n57_w8, 
            w9=> c0_n57_w9, 
            w10=> c0_n57_w10, 
            w11=> c0_n57_w11, 
            w12=> c0_n57_w12, 
            w13=> c0_n57_w13, 
            w14=> c0_n57_w14, 
            w15=> c0_n57_w15, 
            w16=> c0_n57_w16, 
            w17=> c0_n57_w17, 
            w18=> c0_n57_w18, 
            w19=> c0_n57_w19, 
            w20=> c0_n57_w20, 
            w21=> c0_n57_w21, 
            w22=> c0_n57_w22, 
            w23=> c0_n57_w23, 
            w24=> c0_n57_w24, 
            w25=> c0_n57_w25, 
            w26=> c0_n57_w26, 
            w27=> c0_n57_w27, 
            w28=> c0_n57_w28, 
            w29=> c0_n57_w29, 
            w30=> c0_n57_w30, 
            w31=> c0_n57_w31, 
            w32=> c0_n57_w32, 
            w33=> c0_n57_w33, 
            w34=> c0_n57_w34, 
            w35=> c0_n57_w35, 
            w36=> c0_n57_w36, 
            w37=> c0_n57_w37, 
            w38=> c0_n57_w38, 
            w39=> c0_n57_w39, 
            w40=> c0_n57_w40, 
            w41=> c0_n57_w41, 
            w42=> c0_n57_w42, 
            w43=> c0_n57_w43, 
            w44=> c0_n57_w44, 
            w45=> c0_n57_w45, 
            w46=> c0_n57_w46, 
            w47=> c0_n57_w47, 
            w48=> c0_n57_w48, 
            w49=> c0_n57_w49, 
            w50=> c0_n57_w50, 
            w51=> c0_n57_w51, 
            w52=> c0_n57_w52, 
            w53=> c0_n57_w53, 
            w54=> c0_n57_w54, 
            w55=> c0_n57_w55, 
            w56=> c0_n57_w56, 
            w57=> c0_n57_w57, 
            w58=> c0_n57_w58, 
            w59=> c0_n57_w59, 
            w60=> c0_n57_w60, 
            w61=> c0_n57_w61, 
            w62=> c0_n57_w62, 
            w63=> c0_n57_w63, 
            w64=> c0_n57_w64, 
            w65=> c0_n57_w65, 
            w66=> c0_n57_w66, 
            w67=> c0_n57_w67, 
            w68=> c0_n57_w68, 
            w69=> c0_n57_w69, 
            w70=> c0_n57_w70, 
            w71=> c0_n57_w71, 
            w72=> c0_n57_w72, 
            w73=> c0_n57_w73, 
            w74=> c0_n57_w74, 
            w75=> c0_n57_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n57_y
   );           
            
neuron_inst_58: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n58_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n58_w1, 
            w2=> c0_n58_w2, 
            w3=> c0_n58_w3, 
            w4=> c0_n58_w4, 
            w5=> c0_n58_w5, 
            w6=> c0_n58_w6, 
            w7=> c0_n58_w7, 
            w8=> c0_n58_w8, 
            w9=> c0_n58_w9, 
            w10=> c0_n58_w10, 
            w11=> c0_n58_w11, 
            w12=> c0_n58_w12, 
            w13=> c0_n58_w13, 
            w14=> c0_n58_w14, 
            w15=> c0_n58_w15, 
            w16=> c0_n58_w16, 
            w17=> c0_n58_w17, 
            w18=> c0_n58_w18, 
            w19=> c0_n58_w19, 
            w20=> c0_n58_w20, 
            w21=> c0_n58_w21, 
            w22=> c0_n58_w22, 
            w23=> c0_n58_w23, 
            w24=> c0_n58_w24, 
            w25=> c0_n58_w25, 
            w26=> c0_n58_w26, 
            w27=> c0_n58_w27, 
            w28=> c0_n58_w28, 
            w29=> c0_n58_w29, 
            w30=> c0_n58_w30, 
            w31=> c0_n58_w31, 
            w32=> c0_n58_w32, 
            w33=> c0_n58_w33, 
            w34=> c0_n58_w34, 
            w35=> c0_n58_w35, 
            w36=> c0_n58_w36, 
            w37=> c0_n58_w37, 
            w38=> c0_n58_w38, 
            w39=> c0_n58_w39, 
            w40=> c0_n58_w40, 
            w41=> c0_n58_w41, 
            w42=> c0_n58_w42, 
            w43=> c0_n58_w43, 
            w44=> c0_n58_w44, 
            w45=> c0_n58_w45, 
            w46=> c0_n58_w46, 
            w47=> c0_n58_w47, 
            w48=> c0_n58_w48, 
            w49=> c0_n58_w49, 
            w50=> c0_n58_w50, 
            w51=> c0_n58_w51, 
            w52=> c0_n58_w52, 
            w53=> c0_n58_w53, 
            w54=> c0_n58_w54, 
            w55=> c0_n58_w55, 
            w56=> c0_n58_w56, 
            w57=> c0_n58_w57, 
            w58=> c0_n58_w58, 
            w59=> c0_n58_w59, 
            w60=> c0_n58_w60, 
            w61=> c0_n58_w61, 
            w62=> c0_n58_w62, 
            w63=> c0_n58_w63, 
            w64=> c0_n58_w64, 
            w65=> c0_n58_w65, 
            w66=> c0_n58_w66, 
            w67=> c0_n58_w67, 
            w68=> c0_n58_w68, 
            w69=> c0_n58_w69, 
            w70=> c0_n58_w70, 
            w71=> c0_n58_w71, 
            w72=> c0_n58_w72, 
            w73=> c0_n58_w73, 
            w74=> c0_n58_w74, 
            w75=> c0_n58_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n58_y
   );           
            
neuron_inst_59: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n59_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n59_w1, 
            w2=> c0_n59_w2, 
            w3=> c0_n59_w3, 
            w4=> c0_n59_w4, 
            w5=> c0_n59_w5, 
            w6=> c0_n59_w6, 
            w7=> c0_n59_w7, 
            w8=> c0_n59_w8, 
            w9=> c0_n59_w9, 
            w10=> c0_n59_w10, 
            w11=> c0_n59_w11, 
            w12=> c0_n59_w12, 
            w13=> c0_n59_w13, 
            w14=> c0_n59_w14, 
            w15=> c0_n59_w15, 
            w16=> c0_n59_w16, 
            w17=> c0_n59_w17, 
            w18=> c0_n59_w18, 
            w19=> c0_n59_w19, 
            w20=> c0_n59_w20, 
            w21=> c0_n59_w21, 
            w22=> c0_n59_w22, 
            w23=> c0_n59_w23, 
            w24=> c0_n59_w24, 
            w25=> c0_n59_w25, 
            w26=> c0_n59_w26, 
            w27=> c0_n59_w27, 
            w28=> c0_n59_w28, 
            w29=> c0_n59_w29, 
            w30=> c0_n59_w30, 
            w31=> c0_n59_w31, 
            w32=> c0_n59_w32, 
            w33=> c0_n59_w33, 
            w34=> c0_n59_w34, 
            w35=> c0_n59_w35, 
            w36=> c0_n59_w36, 
            w37=> c0_n59_w37, 
            w38=> c0_n59_w38, 
            w39=> c0_n59_w39, 
            w40=> c0_n59_w40, 
            w41=> c0_n59_w41, 
            w42=> c0_n59_w42, 
            w43=> c0_n59_w43, 
            w44=> c0_n59_w44, 
            w45=> c0_n59_w45, 
            w46=> c0_n59_w46, 
            w47=> c0_n59_w47, 
            w48=> c0_n59_w48, 
            w49=> c0_n59_w49, 
            w50=> c0_n59_w50, 
            w51=> c0_n59_w51, 
            w52=> c0_n59_w52, 
            w53=> c0_n59_w53, 
            w54=> c0_n59_w54, 
            w55=> c0_n59_w55, 
            w56=> c0_n59_w56, 
            w57=> c0_n59_w57, 
            w58=> c0_n59_w58, 
            w59=> c0_n59_w59, 
            w60=> c0_n59_w60, 
            w61=> c0_n59_w61, 
            w62=> c0_n59_w62, 
            w63=> c0_n59_w63, 
            w64=> c0_n59_w64, 
            w65=> c0_n59_w65, 
            w66=> c0_n59_w66, 
            w67=> c0_n59_w67, 
            w68=> c0_n59_w68, 
            w69=> c0_n59_w69, 
            w70=> c0_n59_w70, 
            w71=> c0_n59_w71, 
            w72=> c0_n59_w72, 
            w73=> c0_n59_w73, 
            w74=> c0_n59_w74, 
            w75=> c0_n59_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n59_y
   );           
            
neuron_inst_60: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n60_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n60_w1, 
            w2=> c0_n60_w2, 
            w3=> c0_n60_w3, 
            w4=> c0_n60_w4, 
            w5=> c0_n60_w5, 
            w6=> c0_n60_w6, 
            w7=> c0_n60_w7, 
            w8=> c0_n60_w8, 
            w9=> c0_n60_w9, 
            w10=> c0_n60_w10, 
            w11=> c0_n60_w11, 
            w12=> c0_n60_w12, 
            w13=> c0_n60_w13, 
            w14=> c0_n60_w14, 
            w15=> c0_n60_w15, 
            w16=> c0_n60_w16, 
            w17=> c0_n60_w17, 
            w18=> c0_n60_w18, 
            w19=> c0_n60_w19, 
            w20=> c0_n60_w20, 
            w21=> c0_n60_w21, 
            w22=> c0_n60_w22, 
            w23=> c0_n60_w23, 
            w24=> c0_n60_w24, 
            w25=> c0_n60_w25, 
            w26=> c0_n60_w26, 
            w27=> c0_n60_w27, 
            w28=> c0_n60_w28, 
            w29=> c0_n60_w29, 
            w30=> c0_n60_w30, 
            w31=> c0_n60_w31, 
            w32=> c0_n60_w32, 
            w33=> c0_n60_w33, 
            w34=> c0_n60_w34, 
            w35=> c0_n60_w35, 
            w36=> c0_n60_w36, 
            w37=> c0_n60_w37, 
            w38=> c0_n60_w38, 
            w39=> c0_n60_w39, 
            w40=> c0_n60_w40, 
            w41=> c0_n60_w41, 
            w42=> c0_n60_w42, 
            w43=> c0_n60_w43, 
            w44=> c0_n60_w44, 
            w45=> c0_n60_w45, 
            w46=> c0_n60_w46, 
            w47=> c0_n60_w47, 
            w48=> c0_n60_w48, 
            w49=> c0_n60_w49, 
            w50=> c0_n60_w50, 
            w51=> c0_n60_w51, 
            w52=> c0_n60_w52, 
            w53=> c0_n60_w53, 
            w54=> c0_n60_w54, 
            w55=> c0_n60_w55, 
            w56=> c0_n60_w56, 
            w57=> c0_n60_w57, 
            w58=> c0_n60_w58, 
            w59=> c0_n60_w59, 
            w60=> c0_n60_w60, 
            w61=> c0_n60_w61, 
            w62=> c0_n60_w62, 
            w63=> c0_n60_w63, 
            w64=> c0_n60_w64, 
            w65=> c0_n60_w65, 
            w66=> c0_n60_w66, 
            w67=> c0_n60_w67, 
            w68=> c0_n60_w68, 
            w69=> c0_n60_w69, 
            w70=> c0_n60_w70, 
            w71=> c0_n60_w71, 
            w72=> c0_n60_w72, 
            w73=> c0_n60_w73, 
            w74=> c0_n60_w74, 
            w75=> c0_n60_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n60_y
   );           
            
neuron_inst_61: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n61_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n61_w1, 
            w2=> c0_n61_w2, 
            w3=> c0_n61_w3, 
            w4=> c0_n61_w4, 
            w5=> c0_n61_w5, 
            w6=> c0_n61_w6, 
            w7=> c0_n61_w7, 
            w8=> c0_n61_w8, 
            w9=> c0_n61_w9, 
            w10=> c0_n61_w10, 
            w11=> c0_n61_w11, 
            w12=> c0_n61_w12, 
            w13=> c0_n61_w13, 
            w14=> c0_n61_w14, 
            w15=> c0_n61_w15, 
            w16=> c0_n61_w16, 
            w17=> c0_n61_w17, 
            w18=> c0_n61_w18, 
            w19=> c0_n61_w19, 
            w20=> c0_n61_w20, 
            w21=> c0_n61_w21, 
            w22=> c0_n61_w22, 
            w23=> c0_n61_w23, 
            w24=> c0_n61_w24, 
            w25=> c0_n61_w25, 
            w26=> c0_n61_w26, 
            w27=> c0_n61_w27, 
            w28=> c0_n61_w28, 
            w29=> c0_n61_w29, 
            w30=> c0_n61_w30, 
            w31=> c0_n61_w31, 
            w32=> c0_n61_w32, 
            w33=> c0_n61_w33, 
            w34=> c0_n61_w34, 
            w35=> c0_n61_w35, 
            w36=> c0_n61_w36, 
            w37=> c0_n61_w37, 
            w38=> c0_n61_w38, 
            w39=> c0_n61_w39, 
            w40=> c0_n61_w40, 
            w41=> c0_n61_w41, 
            w42=> c0_n61_w42, 
            w43=> c0_n61_w43, 
            w44=> c0_n61_w44, 
            w45=> c0_n61_w45, 
            w46=> c0_n61_w46, 
            w47=> c0_n61_w47, 
            w48=> c0_n61_w48, 
            w49=> c0_n61_w49, 
            w50=> c0_n61_w50, 
            w51=> c0_n61_w51, 
            w52=> c0_n61_w52, 
            w53=> c0_n61_w53, 
            w54=> c0_n61_w54, 
            w55=> c0_n61_w55, 
            w56=> c0_n61_w56, 
            w57=> c0_n61_w57, 
            w58=> c0_n61_w58, 
            w59=> c0_n61_w59, 
            w60=> c0_n61_w60, 
            w61=> c0_n61_w61, 
            w62=> c0_n61_w62, 
            w63=> c0_n61_w63, 
            w64=> c0_n61_w64, 
            w65=> c0_n61_w65, 
            w66=> c0_n61_w66, 
            w67=> c0_n61_w67, 
            w68=> c0_n61_w68, 
            w69=> c0_n61_w69, 
            w70=> c0_n61_w70, 
            w71=> c0_n61_w71, 
            w72=> c0_n61_w72, 
            w73=> c0_n61_w73, 
            w74=> c0_n61_w74, 
            w75=> c0_n61_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n61_y
   );           
            
neuron_inst_62: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n62_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n62_w1, 
            w2=> c0_n62_w2, 
            w3=> c0_n62_w3, 
            w4=> c0_n62_w4, 
            w5=> c0_n62_w5, 
            w6=> c0_n62_w6, 
            w7=> c0_n62_w7, 
            w8=> c0_n62_w8, 
            w9=> c0_n62_w9, 
            w10=> c0_n62_w10, 
            w11=> c0_n62_w11, 
            w12=> c0_n62_w12, 
            w13=> c0_n62_w13, 
            w14=> c0_n62_w14, 
            w15=> c0_n62_w15, 
            w16=> c0_n62_w16, 
            w17=> c0_n62_w17, 
            w18=> c0_n62_w18, 
            w19=> c0_n62_w19, 
            w20=> c0_n62_w20, 
            w21=> c0_n62_w21, 
            w22=> c0_n62_w22, 
            w23=> c0_n62_w23, 
            w24=> c0_n62_w24, 
            w25=> c0_n62_w25, 
            w26=> c0_n62_w26, 
            w27=> c0_n62_w27, 
            w28=> c0_n62_w28, 
            w29=> c0_n62_w29, 
            w30=> c0_n62_w30, 
            w31=> c0_n62_w31, 
            w32=> c0_n62_w32, 
            w33=> c0_n62_w33, 
            w34=> c0_n62_w34, 
            w35=> c0_n62_w35, 
            w36=> c0_n62_w36, 
            w37=> c0_n62_w37, 
            w38=> c0_n62_w38, 
            w39=> c0_n62_w39, 
            w40=> c0_n62_w40, 
            w41=> c0_n62_w41, 
            w42=> c0_n62_w42, 
            w43=> c0_n62_w43, 
            w44=> c0_n62_w44, 
            w45=> c0_n62_w45, 
            w46=> c0_n62_w46, 
            w47=> c0_n62_w47, 
            w48=> c0_n62_w48, 
            w49=> c0_n62_w49, 
            w50=> c0_n62_w50, 
            w51=> c0_n62_w51, 
            w52=> c0_n62_w52, 
            w53=> c0_n62_w53, 
            w54=> c0_n62_w54, 
            w55=> c0_n62_w55, 
            w56=> c0_n62_w56, 
            w57=> c0_n62_w57, 
            w58=> c0_n62_w58, 
            w59=> c0_n62_w59, 
            w60=> c0_n62_w60, 
            w61=> c0_n62_w61, 
            w62=> c0_n62_w62, 
            w63=> c0_n62_w63, 
            w64=> c0_n62_w64, 
            w65=> c0_n62_w65, 
            w66=> c0_n62_w66, 
            w67=> c0_n62_w67, 
            w68=> c0_n62_w68, 
            w69=> c0_n62_w69, 
            w70=> c0_n62_w70, 
            w71=> c0_n62_w71, 
            w72=> c0_n62_w72, 
            w73=> c0_n62_w73, 
            w74=> c0_n62_w74, 
            w75=> c0_n62_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n62_y
   );           
            
neuron_inst_63: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n63_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n63_w1, 
            w2=> c0_n63_w2, 
            w3=> c0_n63_w3, 
            w4=> c0_n63_w4, 
            w5=> c0_n63_w5, 
            w6=> c0_n63_w6, 
            w7=> c0_n63_w7, 
            w8=> c0_n63_w8, 
            w9=> c0_n63_w9, 
            w10=> c0_n63_w10, 
            w11=> c0_n63_w11, 
            w12=> c0_n63_w12, 
            w13=> c0_n63_w13, 
            w14=> c0_n63_w14, 
            w15=> c0_n63_w15, 
            w16=> c0_n63_w16, 
            w17=> c0_n63_w17, 
            w18=> c0_n63_w18, 
            w19=> c0_n63_w19, 
            w20=> c0_n63_w20, 
            w21=> c0_n63_w21, 
            w22=> c0_n63_w22, 
            w23=> c0_n63_w23, 
            w24=> c0_n63_w24, 
            w25=> c0_n63_w25, 
            w26=> c0_n63_w26, 
            w27=> c0_n63_w27, 
            w28=> c0_n63_w28, 
            w29=> c0_n63_w29, 
            w30=> c0_n63_w30, 
            w31=> c0_n63_w31, 
            w32=> c0_n63_w32, 
            w33=> c0_n63_w33, 
            w34=> c0_n63_w34, 
            w35=> c0_n63_w35, 
            w36=> c0_n63_w36, 
            w37=> c0_n63_w37, 
            w38=> c0_n63_w38, 
            w39=> c0_n63_w39, 
            w40=> c0_n63_w40, 
            w41=> c0_n63_w41, 
            w42=> c0_n63_w42, 
            w43=> c0_n63_w43, 
            w44=> c0_n63_w44, 
            w45=> c0_n63_w45, 
            w46=> c0_n63_w46, 
            w47=> c0_n63_w47, 
            w48=> c0_n63_w48, 
            w49=> c0_n63_w49, 
            w50=> c0_n63_w50, 
            w51=> c0_n63_w51, 
            w52=> c0_n63_w52, 
            w53=> c0_n63_w53, 
            w54=> c0_n63_w54, 
            w55=> c0_n63_w55, 
            w56=> c0_n63_w56, 
            w57=> c0_n63_w57, 
            w58=> c0_n63_w58, 
            w59=> c0_n63_w59, 
            w60=> c0_n63_w60, 
            w61=> c0_n63_w61, 
            w62=> c0_n63_w62, 
            w63=> c0_n63_w63, 
            w64=> c0_n63_w64, 
            w65=> c0_n63_w65, 
            w66=> c0_n63_w66, 
            w67=> c0_n63_w67, 
            w68=> c0_n63_w68, 
            w69=> c0_n63_w69, 
            w70=> c0_n63_w70, 
            w71=> c0_n63_w71, 
            w72=> c0_n63_w72, 
            w73=> c0_n63_w73, 
            w74=> c0_n63_w74, 
            w75=> c0_n63_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n63_y
   );           
            
neuron_inst_64: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n64_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n64_w1, 
            w2=> c0_n64_w2, 
            w3=> c0_n64_w3, 
            w4=> c0_n64_w4, 
            w5=> c0_n64_w5, 
            w6=> c0_n64_w6, 
            w7=> c0_n64_w7, 
            w8=> c0_n64_w8, 
            w9=> c0_n64_w9, 
            w10=> c0_n64_w10, 
            w11=> c0_n64_w11, 
            w12=> c0_n64_w12, 
            w13=> c0_n64_w13, 
            w14=> c0_n64_w14, 
            w15=> c0_n64_w15, 
            w16=> c0_n64_w16, 
            w17=> c0_n64_w17, 
            w18=> c0_n64_w18, 
            w19=> c0_n64_w19, 
            w20=> c0_n64_w20, 
            w21=> c0_n64_w21, 
            w22=> c0_n64_w22, 
            w23=> c0_n64_w23, 
            w24=> c0_n64_w24, 
            w25=> c0_n64_w25, 
            w26=> c0_n64_w26, 
            w27=> c0_n64_w27, 
            w28=> c0_n64_w28, 
            w29=> c0_n64_w29, 
            w30=> c0_n64_w30, 
            w31=> c0_n64_w31, 
            w32=> c0_n64_w32, 
            w33=> c0_n64_w33, 
            w34=> c0_n64_w34, 
            w35=> c0_n64_w35, 
            w36=> c0_n64_w36, 
            w37=> c0_n64_w37, 
            w38=> c0_n64_w38, 
            w39=> c0_n64_w39, 
            w40=> c0_n64_w40, 
            w41=> c0_n64_w41, 
            w42=> c0_n64_w42, 
            w43=> c0_n64_w43, 
            w44=> c0_n64_w44, 
            w45=> c0_n64_w45, 
            w46=> c0_n64_w46, 
            w47=> c0_n64_w47, 
            w48=> c0_n64_w48, 
            w49=> c0_n64_w49, 
            w50=> c0_n64_w50, 
            w51=> c0_n64_w51, 
            w52=> c0_n64_w52, 
            w53=> c0_n64_w53, 
            w54=> c0_n64_w54, 
            w55=> c0_n64_w55, 
            w56=> c0_n64_w56, 
            w57=> c0_n64_w57, 
            w58=> c0_n64_w58, 
            w59=> c0_n64_w59, 
            w60=> c0_n64_w60, 
            w61=> c0_n64_w61, 
            w62=> c0_n64_w62, 
            w63=> c0_n64_w63, 
            w64=> c0_n64_w64, 
            w65=> c0_n64_w65, 
            w66=> c0_n64_w66, 
            w67=> c0_n64_w67, 
            w68=> c0_n64_w68, 
            w69=> c0_n64_w69, 
            w70=> c0_n64_w70, 
            w71=> c0_n64_w71, 
            w72=> c0_n64_w72, 
            w73=> c0_n64_w73, 
            w74=> c0_n64_w74, 
            w75=> c0_n64_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n64_y
   );           
            
neuron_inst_65: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n65_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n65_w1, 
            w2=> c0_n65_w2, 
            w3=> c0_n65_w3, 
            w4=> c0_n65_w4, 
            w5=> c0_n65_w5, 
            w6=> c0_n65_w6, 
            w7=> c0_n65_w7, 
            w8=> c0_n65_w8, 
            w9=> c0_n65_w9, 
            w10=> c0_n65_w10, 
            w11=> c0_n65_w11, 
            w12=> c0_n65_w12, 
            w13=> c0_n65_w13, 
            w14=> c0_n65_w14, 
            w15=> c0_n65_w15, 
            w16=> c0_n65_w16, 
            w17=> c0_n65_w17, 
            w18=> c0_n65_w18, 
            w19=> c0_n65_w19, 
            w20=> c0_n65_w20, 
            w21=> c0_n65_w21, 
            w22=> c0_n65_w22, 
            w23=> c0_n65_w23, 
            w24=> c0_n65_w24, 
            w25=> c0_n65_w25, 
            w26=> c0_n65_w26, 
            w27=> c0_n65_w27, 
            w28=> c0_n65_w28, 
            w29=> c0_n65_w29, 
            w30=> c0_n65_w30, 
            w31=> c0_n65_w31, 
            w32=> c0_n65_w32, 
            w33=> c0_n65_w33, 
            w34=> c0_n65_w34, 
            w35=> c0_n65_w35, 
            w36=> c0_n65_w36, 
            w37=> c0_n65_w37, 
            w38=> c0_n65_w38, 
            w39=> c0_n65_w39, 
            w40=> c0_n65_w40, 
            w41=> c0_n65_w41, 
            w42=> c0_n65_w42, 
            w43=> c0_n65_w43, 
            w44=> c0_n65_w44, 
            w45=> c0_n65_w45, 
            w46=> c0_n65_w46, 
            w47=> c0_n65_w47, 
            w48=> c0_n65_w48, 
            w49=> c0_n65_w49, 
            w50=> c0_n65_w50, 
            w51=> c0_n65_w51, 
            w52=> c0_n65_w52, 
            w53=> c0_n65_w53, 
            w54=> c0_n65_w54, 
            w55=> c0_n65_w55, 
            w56=> c0_n65_w56, 
            w57=> c0_n65_w57, 
            w58=> c0_n65_w58, 
            w59=> c0_n65_w59, 
            w60=> c0_n65_w60, 
            w61=> c0_n65_w61, 
            w62=> c0_n65_w62, 
            w63=> c0_n65_w63, 
            w64=> c0_n65_w64, 
            w65=> c0_n65_w65, 
            w66=> c0_n65_w66, 
            w67=> c0_n65_w67, 
            w68=> c0_n65_w68, 
            w69=> c0_n65_w69, 
            w70=> c0_n65_w70, 
            w71=> c0_n65_w71, 
            w72=> c0_n65_w72, 
            w73=> c0_n65_w73, 
            w74=> c0_n65_w74, 
            w75=> c0_n65_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n65_y
   );           
            
neuron_inst_66: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n66_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n66_w1, 
            w2=> c0_n66_w2, 
            w3=> c0_n66_w3, 
            w4=> c0_n66_w4, 
            w5=> c0_n66_w5, 
            w6=> c0_n66_w6, 
            w7=> c0_n66_w7, 
            w8=> c0_n66_w8, 
            w9=> c0_n66_w9, 
            w10=> c0_n66_w10, 
            w11=> c0_n66_w11, 
            w12=> c0_n66_w12, 
            w13=> c0_n66_w13, 
            w14=> c0_n66_w14, 
            w15=> c0_n66_w15, 
            w16=> c0_n66_w16, 
            w17=> c0_n66_w17, 
            w18=> c0_n66_w18, 
            w19=> c0_n66_w19, 
            w20=> c0_n66_w20, 
            w21=> c0_n66_w21, 
            w22=> c0_n66_w22, 
            w23=> c0_n66_w23, 
            w24=> c0_n66_w24, 
            w25=> c0_n66_w25, 
            w26=> c0_n66_w26, 
            w27=> c0_n66_w27, 
            w28=> c0_n66_w28, 
            w29=> c0_n66_w29, 
            w30=> c0_n66_w30, 
            w31=> c0_n66_w31, 
            w32=> c0_n66_w32, 
            w33=> c0_n66_w33, 
            w34=> c0_n66_w34, 
            w35=> c0_n66_w35, 
            w36=> c0_n66_w36, 
            w37=> c0_n66_w37, 
            w38=> c0_n66_w38, 
            w39=> c0_n66_w39, 
            w40=> c0_n66_w40, 
            w41=> c0_n66_w41, 
            w42=> c0_n66_w42, 
            w43=> c0_n66_w43, 
            w44=> c0_n66_w44, 
            w45=> c0_n66_w45, 
            w46=> c0_n66_w46, 
            w47=> c0_n66_w47, 
            w48=> c0_n66_w48, 
            w49=> c0_n66_w49, 
            w50=> c0_n66_w50, 
            w51=> c0_n66_w51, 
            w52=> c0_n66_w52, 
            w53=> c0_n66_w53, 
            w54=> c0_n66_w54, 
            w55=> c0_n66_w55, 
            w56=> c0_n66_w56, 
            w57=> c0_n66_w57, 
            w58=> c0_n66_w58, 
            w59=> c0_n66_w59, 
            w60=> c0_n66_w60, 
            w61=> c0_n66_w61, 
            w62=> c0_n66_w62, 
            w63=> c0_n66_w63, 
            w64=> c0_n66_w64, 
            w65=> c0_n66_w65, 
            w66=> c0_n66_w66, 
            w67=> c0_n66_w67, 
            w68=> c0_n66_w68, 
            w69=> c0_n66_w69, 
            w70=> c0_n66_w70, 
            w71=> c0_n66_w71, 
            w72=> c0_n66_w72, 
            w73=> c0_n66_w73, 
            w74=> c0_n66_w74, 
            w75=> c0_n66_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n66_y
   );           
            
neuron_inst_67: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n67_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n67_w1, 
            w2=> c0_n67_w2, 
            w3=> c0_n67_w3, 
            w4=> c0_n67_w4, 
            w5=> c0_n67_w5, 
            w6=> c0_n67_w6, 
            w7=> c0_n67_w7, 
            w8=> c0_n67_w8, 
            w9=> c0_n67_w9, 
            w10=> c0_n67_w10, 
            w11=> c0_n67_w11, 
            w12=> c0_n67_w12, 
            w13=> c0_n67_w13, 
            w14=> c0_n67_w14, 
            w15=> c0_n67_w15, 
            w16=> c0_n67_w16, 
            w17=> c0_n67_w17, 
            w18=> c0_n67_w18, 
            w19=> c0_n67_w19, 
            w20=> c0_n67_w20, 
            w21=> c0_n67_w21, 
            w22=> c0_n67_w22, 
            w23=> c0_n67_w23, 
            w24=> c0_n67_w24, 
            w25=> c0_n67_w25, 
            w26=> c0_n67_w26, 
            w27=> c0_n67_w27, 
            w28=> c0_n67_w28, 
            w29=> c0_n67_w29, 
            w30=> c0_n67_w30, 
            w31=> c0_n67_w31, 
            w32=> c0_n67_w32, 
            w33=> c0_n67_w33, 
            w34=> c0_n67_w34, 
            w35=> c0_n67_w35, 
            w36=> c0_n67_w36, 
            w37=> c0_n67_w37, 
            w38=> c0_n67_w38, 
            w39=> c0_n67_w39, 
            w40=> c0_n67_w40, 
            w41=> c0_n67_w41, 
            w42=> c0_n67_w42, 
            w43=> c0_n67_w43, 
            w44=> c0_n67_w44, 
            w45=> c0_n67_w45, 
            w46=> c0_n67_w46, 
            w47=> c0_n67_w47, 
            w48=> c0_n67_w48, 
            w49=> c0_n67_w49, 
            w50=> c0_n67_w50, 
            w51=> c0_n67_w51, 
            w52=> c0_n67_w52, 
            w53=> c0_n67_w53, 
            w54=> c0_n67_w54, 
            w55=> c0_n67_w55, 
            w56=> c0_n67_w56, 
            w57=> c0_n67_w57, 
            w58=> c0_n67_w58, 
            w59=> c0_n67_w59, 
            w60=> c0_n67_w60, 
            w61=> c0_n67_w61, 
            w62=> c0_n67_w62, 
            w63=> c0_n67_w63, 
            w64=> c0_n67_w64, 
            w65=> c0_n67_w65, 
            w66=> c0_n67_w66, 
            w67=> c0_n67_w67, 
            w68=> c0_n67_w68, 
            w69=> c0_n67_w69, 
            w70=> c0_n67_w70, 
            w71=> c0_n67_w71, 
            w72=> c0_n67_w72, 
            w73=> c0_n67_w73, 
            w74=> c0_n67_w74, 
            w75=> c0_n67_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n67_y
   );           
            
neuron_inst_68: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n68_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n68_w1, 
            w2=> c0_n68_w2, 
            w3=> c0_n68_w3, 
            w4=> c0_n68_w4, 
            w5=> c0_n68_w5, 
            w6=> c0_n68_w6, 
            w7=> c0_n68_w7, 
            w8=> c0_n68_w8, 
            w9=> c0_n68_w9, 
            w10=> c0_n68_w10, 
            w11=> c0_n68_w11, 
            w12=> c0_n68_w12, 
            w13=> c0_n68_w13, 
            w14=> c0_n68_w14, 
            w15=> c0_n68_w15, 
            w16=> c0_n68_w16, 
            w17=> c0_n68_w17, 
            w18=> c0_n68_w18, 
            w19=> c0_n68_w19, 
            w20=> c0_n68_w20, 
            w21=> c0_n68_w21, 
            w22=> c0_n68_w22, 
            w23=> c0_n68_w23, 
            w24=> c0_n68_w24, 
            w25=> c0_n68_w25, 
            w26=> c0_n68_w26, 
            w27=> c0_n68_w27, 
            w28=> c0_n68_w28, 
            w29=> c0_n68_w29, 
            w30=> c0_n68_w30, 
            w31=> c0_n68_w31, 
            w32=> c0_n68_w32, 
            w33=> c0_n68_w33, 
            w34=> c0_n68_w34, 
            w35=> c0_n68_w35, 
            w36=> c0_n68_w36, 
            w37=> c0_n68_w37, 
            w38=> c0_n68_w38, 
            w39=> c0_n68_w39, 
            w40=> c0_n68_w40, 
            w41=> c0_n68_w41, 
            w42=> c0_n68_w42, 
            w43=> c0_n68_w43, 
            w44=> c0_n68_w44, 
            w45=> c0_n68_w45, 
            w46=> c0_n68_w46, 
            w47=> c0_n68_w47, 
            w48=> c0_n68_w48, 
            w49=> c0_n68_w49, 
            w50=> c0_n68_w50, 
            w51=> c0_n68_w51, 
            w52=> c0_n68_w52, 
            w53=> c0_n68_w53, 
            w54=> c0_n68_w54, 
            w55=> c0_n68_w55, 
            w56=> c0_n68_w56, 
            w57=> c0_n68_w57, 
            w58=> c0_n68_w58, 
            w59=> c0_n68_w59, 
            w60=> c0_n68_w60, 
            w61=> c0_n68_w61, 
            w62=> c0_n68_w62, 
            w63=> c0_n68_w63, 
            w64=> c0_n68_w64, 
            w65=> c0_n68_w65, 
            w66=> c0_n68_w66, 
            w67=> c0_n68_w67, 
            w68=> c0_n68_w68, 
            w69=> c0_n68_w69, 
            w70=> c0_n68_w70, 
            w71=> c0_n68_w71, 
            w72=> c0_n68_w72, 
            w73=> c0_n68_w73, 
            w74=> c0_n68_w74, 
            w75=> c0_n68_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n68_y
   );           
            
neuron_inst_69: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n69_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n69_w1, 
            w2=> c0_n69_w2, 
            w3=> c0_n69_w3, 
            w4=> c0_n69_w4, 
            w5=> c0_n69_w5, 
            w6=> c0_n69_w6, 
            w7=> c0_n69_w7, 
            w8=> c0_n69_w8, 
            w9=> c0_n69_w9, 
            w10=> c0_n69_w10, 
            w11=> c0_n69_w11, 
            w12=> c0_n69_w12, 
            w13=> c0_n69_w13, 
            w14=> c0_n69_w14, 
            w15=> c0_n69_w15, 
            w16=> c0_n69_w16, 
            w17=> c0_n69_w17, 
            w18=> c0_n69_w18, 
            w19=> c0_n69_w19, 
            w20=> c0_n69_w20, 
            w21=> c0_n69_w21, 
            w22=> c0_n69_w22, 
            w23=> c0_n69_w23, 
            w24=> c0_n69_w24, 
            w25=> c0_n69_w25, 
            w26=> c0_n69_w26, 
            w27=> c0_n69_w27, 
            w28=> c0_n69_w28, 
            w29=> c0_n69_w29, 
            w30=> c0_n69_w30, 
            w31=> c0_n69_w31, 
            w32=> c0_n69_w32, 
            w33=> c0_n69_w33, 
            w34=> c0_n69_w34, 
            w35=> c0_n69_w35, 
            w36=> c0_n69_w36, 
            w37=> c0_n69_w37, 
            w38=> c0_n69_w38, 
            w39=> c0_n69_w39, 
            w40=> c0_n69_w40, 
            w41=> c0_n69_w41, 
            w42=> c0_n69_w42, 
            w43=> c0_n69_w43, 
            w44=> c0_n69_w44, 
            w45=> c0_n69_w45, 
            w46=> c0_n69_w46, 
            w47=> c0_n69_w47, 
            w48=> c0_n69_w48, 
            w49=> c0_n69_w49, 
            w50=> c0_n69_w50, 
            w51=> c0_n69_w51, 
            w52=> c0_n69_w52, 
            w53=> c0_n69_w53, 
            w54=> c0_n69_w54, 
            w55=> c0_n69_w55, 
            w56=> c0_n69_w56, 
            w57=> c0_n69_w57, 
            w58=> c0_n69_w58, 
            w59=> c0_n69_w59, 
            w60=> c0_n69_w60, 
            w61=> c0_n69_w61, 
            w62=> c0_n69_w62, 
            w63=> c0_n69_w63, 
            w64=> c0_n69_w64, 
            w65=> c0_n69_w65, 
            w66=> c0_n69_w66, 
            w67=> c0_n69_w67, 
            w68=> c0_n69_w68, 
            w69=> c0_n69_w69, 
            w70=> c0_n69_w70, 
            w71=> c0_n69_w71, 
            w72=> c0_n69_w72, 
            w73=> c0_n69_w73, 
            w74=> c0_n69_w74, 
            w75=> c0_n69_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n69_y
   );           
            
neuron_inst_70: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n70_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n70_w1, 
            w2=> c0_n70_w2, 
            w3=> c0_n70_w3, 
            w4=> c0_n70_w4, 
            w5=> c0_n70_w5, 
            w6=> c0_n70_w6, 
            w7=> c0_n70_w7, 
            w8=> c0_n70_w8, 
            w9=> c0_n70_w9, 
            w10=> c0_n70_w10, 
            w11=> c0_n70_w11, 
            w12=> c0_n70_w12, 
            w13=> c0_n70_w13, 
            w14=> c0_n70_w14, 
            w15=> c0_n70_w15, 
            w16=> c0_n70_w16, 
            w17=> c0_n70_w17, 
            w18=> c0_n70_w18, 
            w19=> c0_n70_w19, 
            w20=> c0_n70_w20, 
            w21=> c0_n70_w21, 
            w22=> c0_n70_w22, 
            w23=> c0_n70_w23, 
            w24=> c0_n70_w24, 
            w25=> c0_n70_w25, 
            w26=> c0_n70_w26, 
            w27=> c0_n70_w27, 
            w28=> c0_n70_w28, 
            w29=> c0_n70_w29, 
            w30=> c0_n70_w30, 
            w31=> c0_n70_w31, 
            w32=> c0_n70_w32, 
            w33=> c0_n70_w33, 
            w34=> c0_n70_w34, 
            w35=> c0_n70_w35, 
            w36=> c0_n70_w36, 
            w37=> c0_n70_w37, 
            w38=> c0_n70_w38, 
            w39=> c0_n70_w39, 
            w40=> c0_n70_w40, 
            w41=> c0_n70_w41, 
            w42=> c0_n70_w42, 
            w43=> c0_n70_w43, 
            w44=> c0_n70_w44, 
            w45=> c0_n70_w45, 
            w46=> c0_n70_w46, 
            w47=> c0_n70_w47, 
            w48=> c0_n70_w48, 
            w49=> c0_n70_w49, 
            w50=> c0_n70_w50, 
            w51=> c0_n70_w51, 
            w52=> c0_n70_w52, 
            w53=> c0_n70_w53, 
            w54=> c0_n70_w54, 
            w55=> c0_n70_w55, 
            w56=> c0_n70_w56, 
            w57=> c0_n70_w57, 
            w58=> c0_n70_w58, 
            w59=> c0_n70_w59, 
            w60=> c0_n70_w60, 
            w61=> c0_n70_w61, 
            w62=> c0_n70_w62, 
            w63=> c0_n70_w63, 
            w64=> c0_n70_w64, 
            w65=> c0_n70_w65, 
            w66=> c0_n70_w66, 
            w67=> c0_n70_w67, 
            w68=> c0_n70_w68, 
            w69=> c0_n70_w69, 
            w70=> c0_n70_w70, 
            w71=> c0_n70_w71, 
            w72=> c0_n70_w72, 
            w73=> c0_n70_w73, 
            w74=> c0_n70_w74, 
            w75=> c0_n70_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n70_y
   );           
            
neuron_inst_71: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n71_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n71_w1, 
            w2=> c0_n71_w2, 
            w3=> c0_n71_w3, 
            w4=> c0_n71_w4, 
            w5=> c0_n71_w5, 
            w6=> c0_n71_w6, 
            w7=> c0_n71_w7, 
            w8=> c0_n71_w8, 
            w9=> c0_n71_w9, 
            w10=> c0_n71_w10, 
            w11=> c0_n71_w11, 
            w12=> c0_n71_w12, 
            w13=> c0_n71_w13, 
            w14=> c0_n71_w14, 
            w15=> c0_n71_w15, 
            w16=> c0_n71_w16, 
            w17=> c0_n71_w17, 
            w18=> c0_n71_w18, 
            w19=> c0_n71_w19, 
            w20=> c0_n71_w20, 
            w21=> c0_n71_w21, 
            w22=> c0_n71_w22, 
            w23=> c0_n71_w23, 
            w24=> c0_n71_w24, 
            w25=> c0_n71_w25, 
            w26=> c0_n71_w26, 
            w27=> c0_n71_w27, 
            w28=> c0_n71_w28, 
            w29=> c0_n71_w29, 
            w30=> c0_n71_w30, 
            w31=> c0_n71_w31, 
            w32=> c0_n71_w32, 
            w33=> c0_n71_w33, 
            w34=> c0_n71_w34, 
            w35=> c0_n71_w35, 
            w36=> c0_n71_w36, 
            w37=> c0_n71_w37, 
            w38=> c0_n71_w38, 
            w39=> c0_n71_w39, 
            w40=> c0_n71_w40, 
            w41=> c0_n71_w41, 
            w42=> c0_n71_w42, 
            w43=> c0_n71_w43, 
            w44=> c0_n71_w44, 
            w45=> c0_n71_w45, 
            w46=> c0_n71_w46, 
            w47=> c0_n71_w47, 
            w48=> c0_n71_w48, 
            w49=> c0_n71_w49, 
            w50=> c0_n71_w50, 
            w51=> c0_n71_w51, 
            w52=> c0_n71_w52, 
            w53=> c0_n71_w53, 
            w54=> c0_n71_w54, 
            w55=> c0_n71_w55, 
            w56=> c0_n71_w56, 
            w57=> c0_n71_w57, 
            w58=> c0_n71_w58, 
            w59=> c0_n71_w59, 
            w60=> c0_n71_w60, 
            w61=> c0_n71_w61, 
            w62=> c0_n71_w62, 
            w63=> c0_n71_w63, 
            w64=> c0_n71_w64, 
            w65=> c0_n71_w65, 
            w66=> c0_n71_w66, 
            w67=> c0_n71_w67, 
            w68=> c0_n71_w68, 
            w69=> c0_n71_w69, 
            w70=> c0_n71_w70, 
            w71=> c0_n71_w71, 
            w72=> c0_n71_w72, 
            w73=> c0_n71_w73, 
            w74=> c0_n71_w74, 
            w75=> c0_n71_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n71_y
   );           
            
neuron_inst_72: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n72_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n72_w1, 
            w2=> c0_n72_w2, 
            w3=> c0_n72_w3, 
            w4=> c0_n72_w4, 
            w5=> c0_n72_w5, 
            w6=> c0_n72_w6, 
            w7=> c0_n72_w7, 
            w8=> c0_n72_w8, 
            w9=> c0_n72_w9, 
            w10=> c0_n72_w10, 
            w11=> c0_n72_w11, 
            w12=> c0_n72_w12, 
            w13=> c0_n72_w13, 
            w14=> c0_n72_w14, 
            w15=> c0_n72_w15, 
            w16=> c0_n72_w16, 
            w17=> c0_n72_w17, 
            w18=> c0_n72_w18, 
            w19=> c0_n72_w19, 
            w20=> c0_n72_w20, 
            w21=> c0_n72_w21, 
            w22=> c0_n72_w22, 
            w23=> c0_n72_w23, 
            w24=> c0_n72_w24, 
            w25=> c0_n72_w25, 
            w26=> c0_n72_w26, 
            w27=> c0_n72_w27, 
            w28=> c0_n72_w28, 
            w29=> c0_n72_w29, 
            w30=> c0_n72_w30, 
            w31=> c0_n72_w31, 
            w32=> c0_n72_w32, 
            w33=> c0_n72_w33, 
            w34=> c0_n72_w34, 
            w35=> c0_n72_w35, 
            w36=> c0_n72_w36, 
            w37=> c0_n72_w37, 
            w38=> c0_n72_w38, 
            w39=> c0_n72_w39, 
            w40=> c0_n72_w40, 
            w41=> c0_n72_w41, 
            w42=> c0_n72_w42, 
            w43=> c0_n72_w43, 
            w44=> c0_n72_w44, 
            w45=> c0_n72_w45, 
            w46=> c0_n72_w46, 
            w47=> c0_n72_w47, 
            w48=> c0_n72_w48, 
            w49=> c0_n72_w49, 
            w50=> c0_n72_w50, 
            w51=> c0_n72_w51, 
            w52=> c0_n72_w52, 
            w53=> c0_n72_w53, 
            w54=> c0_n72_w54, 
            w55=> c0_n72_w55, 
            w56=> c0_n72_w56, 
            w57=> c0_n72_w57, 
            w58=> c0_n72_w58, 
            w59=> c0_n72_w59, 
            w60=> c0_n72_w60, 
            w61=> c0_n72_w61, 
            w62=> c0_n72_w62, 
            w63=> c0_n72_w63, 
            w64=> c0_n72_w64, 
            w65=> c0_n72_w65, 
            w66=> c0_n72_w66, 
            w67=> c0_n72_w67, 
            w68=> c0_n72_w68, 
            w69=> c0_n72_w69, 
            w70=> c0_n72_w70, 
            w71=> c0_n72_w71, 
            w72=> c0_n72_w72, 
            w73=> c0_n72_w73, 
            w74=> c0_n72_w74, 
            w75=> c0_n72_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n72_y
   );           
            
neuron_inst_73: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n73_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n73_w1, 
            w2=> c0_n73_w2, 
            w3=> c0_n73_w3, 
            w4=> c0_n73_w4, 
            w5=> c0_n73_w5, 
            w6=> c0_n73_w6, 
            w7=> c0_n73_w7, 
            w8=> c0_n73_w8, 
            w9=> c0_n73_w9, 
            w10=> c0_n73_w10, 
            w11=> c0_n73_w11, 
            w12=> c0_n73_w12, 
            w13=> c0_n73_w13, 
            w14=> c0_n73_w14, 
            w15=> c0_n73_w15, 
            w16=> c0_n73_w16, 
            w17=> c0_n73_w17, 
            w18=> c0_n73_w18, 
            w19=> c0_n73_w19, 
            w20=> c0_n73_w20, 
            w21=> c0_n73_w21, 
            w22=> c0_n73_w22, 
            w23=> c0_n73_w23, 
            w24=> c0_n73_w24, 
            w25=> c0_n73_w25, 
            w26=> c0_n73_w26, 
            w27=> c0_n73_w27, 
            w28=> c0_n73_w28, 
            w29=> c0_n73_w29, 
            w30=> c0_n73_w30, 
            w31=> c0_n73_w31, 
            w32=> c0_n73_w32, 
            w33=> c0_n73_w33, 
            w34=> c0_n73_w34, 
            w35=> c0_n73_w35, 
            w36=> c0_n73_w36, 
            w37=> c0_n73_w37, 
            w38=> c0_n73_w38, 
            w39=> c0_n73_w39, 
            w40=> c0_n73_w40, 
            w41=> c0_n73_w41, 
            w42=> c0_n73_w42, 
            w43=> c0_n73_w43, 
            w44=> c0_n73_w44, 
            w45=> c0_n73_w45, 
            w46=> c0_n73_w46, 
            w47=> c0_n73_w47, 
            w48=> c0_n73_w48, 
            w49=> c0_n73_w49, 
            w50=> c0_n73_w50, 
            w51=> c0_n73_w51, 
            w52=> c0_n73_w52, 
            w53=> c0_n73_w53, 
            w54=> c0_n73_w54, 
            w55=> c0_n73_w55, 
            w56=> c0_n73_w56, 
            w57=> c0_n73_w57, 
            w58=> c0_n73_w58, 
            w59=> c0_n73_w59, 
            w60=> c0_n73_w60, 
            w61=> c0_n73_w61, 
            w62=> c0_n73_w62, 
            w63=> c0_n73_w63, 
            w64=> c0_n73_w64, 
            w65=> c0_n73_w65, 
            w66=> c0_n73_w66, 
            w67=> c0_n73_w67, 
            w68=> c0_n73_w68, 
            w69=> c0_n73_w69, 
            w70=> c0_n73_w70, 
            w71=> c0_n73_w71, 
            w72=> c0_n73_w72, 
            w73=> c0_n73_w73, 
            w74=> c0_n73_w74, 
            w75=> c0_n73_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n73_y
   );           
            
neuron_inst_74: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n74_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n74_w1, 
            w2=> c0_n74_w2, 
            w3=> c0_n74_w3, 
            w4=> c0_n74_w4, 
            w5=> c0_n74_w5, 
            w6=> c0_n74_w6, 
            w7=> c0_n74_w7, 
            w8=> c0_n74_w8, 
            w9=> c0_n74_w9, 
            w10=> c0_n74_w10, 
            w11=> c0_n74_w11, 
            w12=> c0_n74_w12, 
            w13=> c0_n74_w13, 
            w14=> c0_n74_w14, 
            w15=> c0_n74_w15, 
            w16=> c0_n74_w16, 
            w17=> c0_n74_w17, 
            w18=> c0_n74_w18, 
            w19=> c0_n74_w19, 
            w20=> c0_n74_w20, 
            w21=> c0_n74_w21, 
            w22=> c0_n74_w22, 
            w23=> c0_n74_w23, 
            w24=> c0_n74_w24, 
            w25=> c0_n74_w25, 
            w26=> c0_n74_w26, 
            w27=> c0_n74_w27, 
            w28=> c0_n74_w28, 
            w29=> c0_n74_w29, 
            w30=> c0_n74_w30, 
            w31=> c0_n74_w31, 
            w32=> c0_n74_w32, 
            w33=> c0_n74_w33, 
            w34=> c0_n74_w34, 
            w35=> c0_n74_w35, 
            w36=> c0_n74_w36, 
            w37=> c0_n74_w37, 
            w38=> c0_n74_w38, 
            w39=> c0_n74_w39, 
            w40=> c0_n74_w40, 
            w41=> c0_n74_w41, 
            w42=> c0_n74_w42, 
            w43=> c0_n74_w43, 
            w44=> c0_n74_w44, 
            w45=> c0_n74_w45, 
            w46=> c0_n74_w46, 
            w47=> c0_n74_w47, 
            w48=> c0_n74_w48, 
            w49=> c0_n74_w49, 
            w50=> c0_n74_w50, 
            w51=> c0_n74_w51, 
            w52=> c0_n74_w52, 
            w53=> c0_n74_w53, 
            w54=> c0_n74_w54, 
            w55=> c0_n74_w55, 
            w56=> c0_n74_w56, 
            w57=> c0_n74_w57, 
            w58=> c0_n74_w58, 
            w59=> c0_n74_w59, 
            w60=> c0_n74_w60, 
            w61=> c0_n74_w61, 
            w62=> c0_n74_w62, 
            w63=> c0_n74_w63, 
            w64=> c0_n74_w64, 
            w65=> c0_n74_w65, 
            w66=> c0_n74_w66, 
            w67=> c0_n74_w67, 
            w68=> c0_n74_w68, 
            w69=> c0_n74_w69, 
            w70=> c0_n74_w70, 
            w71=> c0_n74_w71, 
            w72=> c0_n74_w72, 
            w73=> c0_n74_w73, 
            w74=> c0_n74_w74, 
            w75=> c0_n74_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n74_y
   );           
            
neuron_inst_75: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n75_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n75_w1, 
            w2=> c0_n75_w2, 
            w3=> c0_n75_w3, 
            w4=> c0_n75_w4, 
            w5=> c0_n75_w5, 
            w6=> c0_n75_w6, 
            w7=> c0_n75_w7, 
            w8=> c0_n75_w8, 
            w9=> c0_n75_w9, 
            w10=> c0_n75_w10, 
            w11=> c0_n75_w11, 
            w12=> c0_n75_w12, 
            w13=> c0_n75_w13, 
            w14=> c0_n75_w14, 
            w15=> c0_n75_w15, 
            w16=> c0_n75_w16, 
            w17=> c0_n75_w17, 
            w18=> c0_n75_w18, 
            w19=> c0_n75_w19, 
            w20=> c0_n75_w20, 
            w21=> c0_n75_w21, 
            w22=> c0_n75_w22, 
            w23=> c0_n75_w23, 
            w24=> c0_n75_w24, 
            w25=> c0_n75_w25, 
            w26=> c0_n75_w26, 
            w27=> c0_n75_w27, 
            w28=> c0_n75_w28, 
            w29=> c0_n75_w29, 
            w30=> c0_n75_w30, 
            w31=> c0_n75_w31, 
            w32=> c0_n75_w32, 
            w33=> c0_n75_w33, 
            w34=> c0_n75_w34, 
            w35=> c0_n75_w35, 
            w36=> c0_n75_w36, 
            w37=> c0_n75_w37, 
            w38=> c0_n75_w38, 
            w39=> c0_n75_w39, 
            w40=> c0_n75_w40, 
            w41=> c0_n75_w41, 
            w42=> c0_n75_w42, 
            w43=> c0_n75_w43, 
            w44=> c0_n75_w44, 
            w45=> c0_n75_w45, 
            w46=> c0_n75_w46, 
            w47=> c0_n75_w47, 
            w48=> c0_n75_w48, 
            w49=> c0_n75_w49, 
            w50=> c0_n75_w50, 
            w51=> c0_n75_w51, 
            w52=> c0_n75_w52, 
            w53=> c0_n75_w53, 
            w54=> c0_n75_w54, 
            w55=> c0_n75_w55, 
            w56=> c0_n75_w56, 
            w57=> c0_n75_w57, 
            w58=> c0_n75_w58, 
            w59=> c0_n75_w59, 
            w60=> c0_n75_w60, 
            w61=> c0_n75_w61, 
            w62=> c0_n75_w62, 
            w63=> c0_n75_w63, 
            w64=> c0_n75_w64, 
            w65=> c0_n75_w65, 
            w66=> c0_n75_w66, 
            w67=> c0_n75_w67, 
            w68=> c0_n75_w68, 
            w69=> c0_n75_w69, 
            w70=> c0_n75_w70, 
            w71=> c0_n75_w71, 
            w72=> c0_n75_w72, 
            w73=> c0_n75_w73, 
            w74=> c0_n75_w74, 
            w75=> c0_n75_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n75_y
   );           
            
neuron_inst_76: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n76_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n76_w1, 
            w2=> c0_n76_w2, 
            w3=> c0_n76_w3, 
            w4=> c0_n76_w4, 
            w5=> c0_n76_w5, 
            w6=> c0_n76_w6, 
            w7=> c0_n76_w7, 
            w8=> c0_n76_w8, 
            w9=> c0_n76_w9, 
            w10=> c0_n76_w10, 
            w11=> c0_n76_w11, 
            w12=> c0_n76_w12, 
            w13=> c0_n76_w13, 
            w14=> c0_n76_w14, 
            w15=> c0_n76_w15, 
            w16=> c0_n76_w16, 
            w17=> c0_n76_w17, 
            w18=> c0_n76_w18, 
            w19=> c0_n76_w19, 
            w20=> c0_n76_w20, 
            w21=> c0_n76_w21, 
            w22=> c0_n76_w22, 
            w23=> c0_n76_w23, 
            w24=> c0_n76_w24, 
            w25=> c0_n76_w25, 
            w26=> c0_n76_w26, 
            w27=> c0_n76_w27, 
            w28=> c0_n76_w28, 
            w29=> c0_n76_w29, 
            w30=> c0_n76_w30, 
            w31=> c0_n76_w31, 
            w32=> c0_n76_w32, 
            w33=> c0_n76_w33, 
            w34=> c0_n76_w34, 
            w35=> c0_n76_w35, 
            w36=> c0_n76_w36, 
            w37=> c0_n76_w37, 
            w38=> c0_n76_w38, 
            w39=> c0_n76_w39, 
            w40=> c0_n76_w40, 
            w41=> c0_n76_w41, 
            w42=> c0_n76_w42, 
            w43=> c0_n76_w43, 
            w44=> c0_n76_w44, 
            w45=> c0_n76_w45, 
            w46=> c0_n76_w46, 
            w47=> c0_n76_w47, 
            w48=> c0_n76_w48, 
            w49=> c0_n76_w49, 
            w50=> c0_n76_w50, 
            w51=> c0_n76_w51, 
            w52=> c0_n76_w52, 
            w53=> c0_n76_w53, 
            w54=> c0_n76_w54, 
            w55=> c0_n76_w55, 
            w56=> c0_n76_w56, 
            w57=> c0_n76_w57, 
            w58=> c0_n76_w58, 
            w59=> c0_n76_w59, 
            w60=> c0_n76_w60, 
            w61=> c0_n76_w61, 
            w62=> c0_n76_w62, 
            w63=> c0_n76_w63, 
            w64=> c0_n76_w64, 
            w65=> c0_n76_w65, 
            w66=> c0_n76_w66, 
            w67=> c0_n76_w67, 
            w68=> c0_n76_w68, 
            w69=> c0_n76_w69, 
            w70=> c0_n76_w70, 
            w71=> c0_n76_w71, 
            w72=> c0_n76_w72, 
            w73=> c0_n76_w73, 
            w74=> c0_n76_w74, 
            w75=> c0_n76_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n76_y
   );           
            
neuron_inst_77: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n77_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n77_w1, 
            w2=> c0_n77_w2, 
            w3=> c0_n77_w3, 
            w4=> c0_n77_w4, 
            w5=> c0_n77_w5, 
            w6=> c0_n77_w6, 
            w7=> c0_n77_w7, 
            w8=> c0_n77_w8, 
            w9=> c0_n77_w9, 
            w10=> c0_n77_w10, 
            w11=> c0_n77_w11, 
            w12=> c0_n77_w12, 
            w13=> c0_n77_w13, 
            w14=> c0_n77_w14, 
            w15=> c0_n77_w15, 
            w16=> c0_n77_w16, 
            w17=> c0_n77_w17, 
            w18=> c0_n77_w18, 
            w19=> c0_n77_w19, 
            w20=> c0_n77_w20, 
            w21=> c0_n77_w21, 
            w22=> c0_n77_w22, 
            w23=> c0_n77_w23, 
            w24=> c0_n77_w24, 
            w25=> c0_n77_w25, 
            w26=> c0_n77_w26, 
            w27=> c0_n77_w27, 
            w28=> c0_n77_w28, 
            w29=> c0_n77_w29, 
            w30=> c0_n77_w30, 
            w31=> c0_n77_w31, 
            w32=> c0_n77_w32, 
            w33=> c0_n77_w33, 
            w34=> c0_n77_w34, 
            w35=> c0_n77_w35, 
            w36=> c0_n77_w36, 
            w37=> c0_n77_w37, 
            w38=> c0_n77_w38, 
            w39=> c0_n77_w39, 
            w40=> c0_n77_w40, 
            w41=> c0_n77_w41, 
            w42=> c0_n77_w42, 
            w43=> c0_n77_w43, 
            w44=> c0_n77_w44, 
            w45=> c0_n77_w45, 
            w46=> c0_n77_w46, 
            w47=> c0_n77_w47, 
            w48=> c0_n77_w48, 
            w49=> c0_n77_w49, 
            w50=> c0_n77_w50, 
            w51=> c0_n77_w51, 
            w52=> c0_n77_w52, 
            w53=> c0_n77_w53, 
            w54=> c0_n77_w54, 
            w55=> c0_n77_w55, 
            w56=> c0_n77_w56, 
            w57=> c0_n77_w57, 
            w58=> c0_n77_w58, 
            w59=> c0_n77_w59, 
            w60=> c0_n77_w60, 
            w61=> c0_n77_w61, 
            w62=> c0_n77_w62, 
            w63=> c0_n77_w63, 
            w64=> c0_n77_w64, 
            w65=> c0_n77_w65, 
            w66=> c0_n77_w66, 
            w67=> c0_n77_w67, 
            w68=> c0_n77_w68, 
            w69=> c0_n77_w69, 
            w70=> c0_n77_w70, 
            w71=> c0_n77_w71, 
            w72=> c0_n77_w72, 
            w73=> c0_n77_w73, 
            w74=> c0_n77_w74, 
            w75=> c0_n77_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n77_y
   );           
            
neuron_inst_78: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n78_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n78_w1, 
            w2=> c0_n78_w2, 
            w3=> c0_n78_w3, 
            w4=> c0_n78_w4, 
            w5=> c0_n78_w5, 
            w6=> c0_n78_w6, 
            w7=> c0_n78_w7, 
            w8=> c0_n78_w8, 
            w9=> c0_n78_w9, 
            w10=> c0_n78_w10, 
            w11=> c0_n78_w11, 
            w12=> c0_n78_w12, 
            w13=> c0_n78_w13, 
            w14=> c0_n78_w14, 
            w15=> c0_n78_w15, 
            w16=> c0_n78_w16, 
            w17=> c0_n78_w17, 
            w18=> c0_n78_w18, 
            w19=> c0_n78_w19, 
            w20=> c0_n78_w20, 
            w21=> c0_n78_w21, 
            w22=> c0_n78_w22, 
            w23=> c0_n78_w23, 
            w24=> c0_n78_w24, 
            w25=> c0_n78_w25, 
            w26=> c0_n78_w26, 
            w27=> c0_n78_w27, 
            w28=> c0_n78_w28, 
            w29=> c0_n78_w29, 
            w30=> c0_n78_w30, 
            w31=> c0_n78_w31, 
            w32=> c0_n78_w32, 
            w33=> c0_n78_w33, 
            w34=> c0_n78_w34, 
            w35=> c0_n78_w35, 
            w36=> c0_n78_w36, 
            w37=> c0_n78_w37, 
            w38=> c0_n78_w38, 
            w39=> c0_n78_w39, 
            w40=> c0_n78_w40, 
            w41=> c0_n78_w41, 
            w42=> c0_n78_w42, 
            w43=> c0_n78_w43, 
            w44=> c0_n78_w44, 
            w45=> c0_n78_w45, 
            w46=> c0_n78_w46, 
            w47=> c0_n78_w47, 
            w48=> c0_n78_w48, 
            w49=> c0_n78_w49, 
            w50=> c0_n78_w50, 
            w51=> c0_n78_w51, 
            w52=> c0_n78_w52, 
            w53=> c0_n78_w53, 
            w54=> c0_n78_w54, 
            w55=> c0_n78_w55, 
            w56=> c0_n78_w56, 
            w57=> c0_n78_w57, 
            w58=> c0_n78_w58, 
            w59=> c0_n78_w59, 
            w60=> c0_n78_w60, 
            w61=> c0_n78_w61, 
            w62=> c0_n78_w62, 
            w63=> c0_n78_w63, 
            w64=> c0_n78_w64, 
            w65=> c0_n78_w65, 
            w66=> c0_n78_w66, 
            w67=> c0_n78_w67, 
            w68=> c0_n78_w68, 
            w69=> c0_n78_w69, 
            w70=> c0_n78_w70, 
            w71=> c0_n78_w71, 
            w72=> c0_n78_w72, 
            w73=> c0_n78_w73, 
            w74=> c0_n78_w74, 
            w75=> c0_n78_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n78_y
   );           
            
neuron_inst_79: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n79_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n79_w1, 
            w2=> c0_n79_w2, 
            w3=> c0_n79_w3, 
            w4=> c0_n79_w4, 
            w5=> c0_n79_w5, 
            w6=> c0_n79_w6, 
            w7=> c0_n79_w7, 
            w8=> c0_n79_w8, 
            w9=> c0_n79_w9, 
            w10=> c0_n79_w10, 
            w11=> c0_n79_w11, 
            w12=> c0_n79_w12, 
            w13=> c0_n79_w13, 
            w14=> c0_n79_w14, 
            w15=> c0_n79_w15, 
            w16=> c0_n79_w16, 
            w17=> c0_n79_w17, 
            w18=> c0_n79_w18, 
            w19=> c0_n79_w19, 
            w20=> c0_n79_w20, 
            w21=> c0_n79_w21, 
            w22=> c0_n79_w22, 
            w23=> c0_n79_w23, 
            w24=> c0_n79_w24, 
            w25=> c0_n79_w25, 
            w26=> c0_n79_w26, 
            w27=> c0_n79_w27, 
            w28=> c0_n79_w28, 
            w29=> c0_n79_w29, 
            w30=> c0_n79_w30, 
            w31=> c0_n79_w31, 
            w32=> c0_n79_w32, 
            w33=> c0_n79_w33, 
            w34=> c0_n79_w34, 
            w35=> c0_n79_w35, 
            w36=> c0_n79_w36, 
            w37=> c0_n79_w37, 
            w38=> c0_n79_w38, 
            w39=> c0_n79_w39, 
            w40=> c0_n79_w40, 
            w41=> c0_n79_w41, 
            w42=> c0_n79_w42, 
            w43=> c0_n79_w43, 
            w44=> c0_n79_w44, 
            w45=> c0_n79_w45, 
            w46=> c0_n79_w46, 
            w47=> c0_n79_w47, 
            w48=> c0_n79_w48, 
            w49=> c0_n79_w49, 
            w50=> c0_n79_w50, 
            w51=> c0_n79_w51, 
            w52=> c0_n79_w52, 
            w53=> c0_n79_w53, 
            w54=> c0_n79_w54, 
            w55=> c0_n79_w55, 
            w56=> c0_n79_w56, 
            w57=> c0_n79_w57, 
            w58=> c0_n79_w58, 
            w59=> c0_n79_w59, 
            w60=> c0_n79_w60, 
            w61=> c0_n79_w61, 
            w62=> c0_n79_w62, 
            w63=> c0_n79_w63, 
            w64=> c0_n79_w64, 
            w65=> c0_n79_w65, 
            w66=> c0_n79_w66, 
            w67=> c0_n79_w67, 
            w68=> c0_n79_w68, 
            w69=> c0_n79_w69, 
            w70=> c0_n79_w70, 
            w71=> c0_n79_w71, 
            w72=> c0_n79_w72, 
            w73=> c0_n79_w73, 
            w74=> c0_n79_w74, 
            w75=> c0_n79_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n79_y
   );           
            
neuron_inst_80: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n80_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n80_w1, 
            w2=> c0_n80_w2, 
            w3=> c0_n80_w3, 
            w4=> c0_n80_w4, 
            w5=> c0_n80_w5, 
            w6=> c0_n80_w6, 
            w7=> c0_n80_w7, 
            w8=> c0_n80_w8, 
            w9=> c0_n80_w9, 
            w10=> c0_n80_w10, 
            w11=> c0_n80_w11, 
            w12=> c0_n80_w12, 
            w13=> c0_n80_w13, 
            w14=> c0_n80_w14, 
            w15=> c0_n80_w15, 
            w16=> c0_n80_w16, 
            w17=> c0_n80_w17, 
            w18=> c0_n80_w18, 
            w19=> c0_n80_w19, 
            w20=> c0_n80_w20, 
            w21=> c0_n80_w21, 
            w22=> c0_n80_w22, 
            w23=> c0_n80_w23, 
            w24=> c0_n80_w24, 
            w25=> c0_n80_w25, 
            w26=> c0_n80_w26, 
            w27=> c0_n80_w27, 
            w28=> c0_n80_w28, 
            w29=> c0_n80_w29, 
            w30=> c0_n80_w30, 
            w31=> c0_n80_w31, 
            w32=> c0_n80_w32, 
            w33=> c0_n80_w33, 
            w34=> c0_n80_w34, 
            w35=> c0_n80_w35, 
            w36=> c0_n80_w36, 
            w37=> c0_n80_w37, 
            w38=> c0_n80_w38, 
            w39=> c0_n80_w39, 
            w40=> c0_n80_w40, 
            w41=> c0_n80_w41, 
            w42=> c0_n80_w42, 
            w43=> c0_n80_w43, 
            w44=> c0_n80_w44, 
            w45=> c0_n80_w45, 
            w46=> c0_n80_w46, 
            w47=> c0_n80_w47, 
            w48=> c0_n80_w48, 
            w49=> c0_n80_w49, 
            w50=> c0_n80_w50, 
            w51=> c0_n80_w51, 
            w52=> c0_n80_w52, 
            w53=> c0_n80_w53, 
            w54=> c0_n80_w54, 
            w55=> c0_n80_w55, 
            w56=> c0_n80_w56, 
            w57=> c0_n80_w57, 
            w58=> c0_n80_w58, 
            w59=> c0_n80_w59, 
            w60=> c0_n80_w60, 
            w61=> c0_n80_w61, 
            w62=> c0_n80_w62, 
            w63=> c0_n80_w63, 
            w64=> c0_n80_w64, 
            w65=> c0_n80_w65, 
            w66=> c0_n80_w66, 
            w67=> c0_n80_w67, 
            w68=> c0_n80_w68, 
            w69=> c0_n80_w69, 
            w70=> c0_n80_w70, 
            w71=> c0_n80_w71, 
            w72=> c0_n80_w72, 
            w73=> c0_n80_w73, 
            w74=> c0_n80_w74, 
            w75=> c0_n80_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n80_y
   );           
            
neuron_inst_81: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n81_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n81_w1, 
            w2=> c0_n81_w2, 
            w3=> c0_n81_w3, 
            w4=> c0_n81_w4, 
            w5=> c0_n81_w5, 
            w6=> c0_n81_w6, 
            w7=> c0_n81_w7, 
            w8=> c0_n81_w8, 
            w9=> c0_n81_w9, 
            w10=> c0_n81_w10, 
            w11=> c0_n81_w11, 
            w12=> c0_n81_w12, 
            w13=> c0_n81_w13, 
            w14=> c0_n81_w14, 
            w15=> c0_n81_w15, 
            w16=> c0_n81_w16, 
            w17=> c0_n81_w17, 
            w18=> c0_n81_w18, 
            w19=> c0_n81_w19, 
            w20=> c0_n81_w20, 
            w21=> c0_n81_w21, 
            w22=> c0_n81_w22, 
            w23=> c0_n81_w23, 
            w24=> c0_n81_w24, 
            w25=> c0_n81_w25, 
            w26=> c0_n81_w26, 
            w27=> c0_n81_w27, 
            w28=> c0_n81_w28, 
            w29=> c0_n81_w29, 
            w30=> c0_n81_w30, 
            w31=> c0_n81_w31, 
            w32=> c0_n81_w32, 
            w33=> c0_n81_w33, 
            w34=> c0_n81_w34, 
            w35=> c0_n81_w35, 
            w36=> c0_n81_w36, 
            w37=> c0_n81_w37, 
            w38=> c0_n81_w38, 
            w39=> c0_n81_w39, 
            w40=> c0_n81_w40, 
            w41=> c0_n81_w41, 
            w42=> c0_n81_w42, 
            w43=> c0_n81_w43, 
            w44=> c0_n81_w44, 
            w45=> c0_n81_w45, 
            w46=> c0_n81_w46, 
            w47=> c0_n81_w47, 
            w48=> c0_n81_w48, 
            w49=> c0_n81_w49, 
            w50=> c0_n81_w50, 
            w51=> c0_n81_w51, 
            w52=> c0_n81_w52, 
            w53=> c0_n81_w53, 
            w54=> c0_n81_w54, 
            w55=> c0_n81_w55, 
            w56=> c0_n81_w56, 
            w57=> c0_n81_w57, 
            w58=> c0_n81_w58, 
            w59=> c0_n81_w59, 
            w60=> c0_n81_w60, 
            w61=> c0_n81_w61, 
            w62=> c0_n81_w62, 
            w63=> c0_n81_w63, 
            w64=> c0_n81_w64, 
            w65=> c0_n81_w65, 
            w66=> c0_n81_w66, 
            w67=> c0_n81_w67, 
            w68=> c0_n81_w68, 
            w69=> c0_n81_w69, 
            w70=> c0_n81_w70, 
            w71=> c0_n81_w71, 
            w72=> c0_n81_w72, 
            w73=> c0_n81_w73, 
            w74=> c0_n81_w74, 
            w75=> c0_n81_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n81_y
   );           
            
neuron_inst_82: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n82_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n82_w1, 
            w2=> c0_n82_w2, 
            w3=> c0_n82_w3, 
            w4=> c0_n82_w4, 
            w5=> c0_n82_w5, 
            w6=> c0_n82_w6, 
            w7=> c0_n82_w7, 
            w8=> c0_n82_w8, 
            w9=> c0_n82_w9, 
            w10=> c0_n82_w10, 
            w11=> c0_n82_w11, 
            w12=> c0_n82_w12, 
            w13=> c0_n82_w13, 
            w14=> c0_n82_w14, 
            w15=> c0_n82_w15, 
            w16=> c0_n82_w16, 
            w17=> c0_n82_w17, 
            w18=> c0_n82_w18, 
            w19=> c0_n82_w19, 
            w20=> c0_n82_w20, 
            w21=> c0_n82_w21, 
            w22=> c0_n82_w22, 
            w23=> c0_n82_w23, 
            w24=> c0_n82_w24, 
            w25=> c0_n82_w25, 
            w26=> c0_n82_w26, 
            w27=> c0_n82_w27, 
            w28=> c0_n82_w28, 
            w29=> c0_n82_w29, 
            w30=> c0_n82_w30, 
            w31=> c0_n82_w31, 
            w32=> c0_n82_w32, 
            w33=> c0_n82_w33, 
            w34=> c0_n82_w34, 
            w35=> c0_n82_w35, 
            w36=> c0_n82_w36, 
            w37=> c0_n82_w37, 
            w38=> c0_n82_w38, 
            w39=> c0_n82_w39, 
            w40=> c0_n82_w40, 
            w41=> c0_n82_w41, 
            w42=> c0_n82_w42, 
            w43=> c0_n82_w43, 
            w44=> c0_n82_w44, 
            w45=> c0_n82_w45, 
            w46=> c0_n82_w46, 
            w47=> c0_n82_w47, 
            w48=> c0_n82_w48, 
            w49=> c0_n82_w49, 
            w50=> c0_n82_w50, 
            w51=> c0_n82_w51, 
            w52=> c0_n82_w52, 
            w53=> c0_n82_w53, 
            w54=> c0_n82_w54, 
            w55=> c0_n82_w55, 
            w56=> c0_n82_w56, 
            w57=> c0_n82_w57, 
            w58=> c0_n82_w58, 
            w59=> c0_n82_w59, 
            w60=> c0_n82_w60, 
            w61=> c0_n82_w61, 
            w62=> c0_n82_w62, 
            w63=> c0_n82_w63, 
            w64=> c0_n82_w64, 
            w65=> c0_n82_w65, 
            w66=> c0_n82_w66, 
            w67=> c0_n82_w67, 
            w68=> c0_n82_w68, 
            w69=> c0_n82_w69, 
            w70=> c0_n82_w70, 
            w71=> c0_n82_w71, 
            w72=> c0_n82_w72, 
            w73=> c0_n82_w73, 
            w74=> c0_n82_w74, 
            w75=> c0_n82_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n82_y
   );           
            
neuron_inst_83: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n83_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n83_w1, 
            w2=> c0_n83_w2, 
            w3=> c0_n83_w3, 
            w4=> c0_n83_w4, 
            w5=> c0_n83_w5, 
            w6=> c0_n83_w6, 
            w7=> c0_n83_w7, 
            w8=> c0_n83_w8, 
            w9=> c0_n83_w9, 
            w10=> c0_n83_w10, 
            w11=> c0_n83_w11, 
            w12=> c0_n83_w12, 
            w13=> c0_n83_w13, 
            w14=> c0_n83_w14, 
            w15=> c0_n83_w15, 
            w16=> c0_n83_w16, 
            w17=> c0_n83_w17, 
            w18=> c0_n83_w18, 
            w19=> c0_n83_w19, 
            w20=> c0_n83_w20, 
            w21=> c0_n83_w21, 
            w22=> c0_n83_w22, 
            w23=> c0_n83_w23, 
            w24=> c0_n83_w24, 
            w25=> c0_n83_w25, 
            w26=> c0_n83_w26, 
            w27=> c0_n83_w27, 
            w28=> c0_n83_w28, 
            w29=> c0_n83_w29, 
            w30=> c0_n83_w30, 
            w31=> c0_n83_w31, 
            w32=> c0_n83_w32, 
            w33=> c0_n83_w33, 
            w34=> c0_n83_w34, 
            w35=> c0_n83_w35, 
            w36=> c0_n83_w36, 
            w37=> c0_n83_w37, 
            w38=> c0_n83_w38, 
            w39=> c0_n83_w39, 
            w40=> c0_n83_w40, 
            w41=> c0_n83_w41, 
            w42=> c0_n83_w42, 
            w43=> c0_n83_w43, 
            w44=> c0_n83_w44, 
            w45=> c0_n83_w45, 
            w46=> c0_n83_w46, 
            w47=> c0_n83_w47, 
            w48=> c0_n83_w48, 
            w49=> c0_n83_w49, 
            w50=> c0_n83_w50, 
            w51=> c0_n83_w51, 
            w52=> c0_n83_w52, 
            w53=> c0_n83_w53, 
            w54=> c0_n83_w54, 
            w55=> c0_n83_w55, 
            w56=> c0_n83_w56, 
            w57=> c0_n83_w57, 
            w58=> c0_n83_w58, 
            w59=> c0_n83_w59, 
            w60=> c0_n83_w60, 
            w61=> c0_n83_w61, 
            w62=> c0_n83_w62, 
            w63=> c0_n83_w63, 
            w64=> c0_n83_w64, 
            w65=> c0_n83_w65, 
            w66=> c0_n83_w66, 
            w67=> c0_n83_w67, 
            w68=> c0_n83_w68, 
            w69=> c0_n83_w69, 
            w70=> c0_n83_w70, 
            w71=> c0_n83_w71, 
            w72=> c0_n83_w72, 
            w73=> c0_n83_w73, 
            w74=> c0_n83_w74, 
            w75=> c0_n83_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n83_y
   );           
            
neuron_inst_84: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n84_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n84_w1, 
            w2=> c0_n84_w2, 
            w3=> c0_n84_w3, 
            w4=> c0_n84_w4, 
            w5=> c0_n84_w5, 
            w6=> c0_n84_w6, 
            w7=> c0_n84_w7, 
            w8=> c0_n84_w8, 
            w9=> c0_n84_w9, 
            w10=> c0_n84_w10, 
            w11=> c0_n84_w11, 
            w12=> c0_n84_w12, 
            w13=> c0_n84_w13, 
            w14=> c0_n84_w14, 
            w15=> c0_n84_w15, 
            w16=> c0_n84_w16, 
            w17=> c0_n84_w17, 
            w18=> c0_n84_w18, 
            w19=> c0_n84_w19, 
            w20=> c0_n84_w20, 
            w21=> c0_n84_w21, 
            w22=> c0_n84_w22, 
            w23=> c0_n84_w23, 
            w24=> c0_n84_w24, 
            w25=> c0_n84_w25, 
            w26=> c0_n84_w26, 
            w27=> c0_n84_w27, 
            w28=> c0_n84_w28, 
            w29=> c0_n84_w29, 
            w30=> c0_n84_w30, 
            w31=> c0_n84_w31, 
            w32=> c0_n84_w32, 
            w33=> c0_n84_w33, 
            w34=> c0_n84_w34, 
            w35=> c0_n84_w35, 
            w36=> c0_n84_w36, 
            w37=> c0_n84_w37, 
            w38=> c0_n84_w38, 
            w39=> c0_n84_w39, 
            w40=> c0_n84_w40, 
            w41=> c0_n84_w41, 
            w42=> c0_n84_w42, 
            w43=> c0_n84_w43, 
            w44=> c0_n84_w44, 
            w45=> c0_n84_w45, 
            w46=> c0_n84_w46, 
            w47=> c0_n84_w47, 
            w48=> c0_n84_w48, 
            w49=> c0_n84_w49, 
            w50=> c0_n84_w50, 
            w51=> c0_n84_w51, 
            w52=> c0_n84_w52, 
            w53=> c0_n84_w53, 
            w54=> c0_n84_w54, 
            w55=> c0_n84_w55, 
            w56=> c0_n84_w56, 
            w57=> c0_n84_w57, 
            w58=> c0_n84_w58, 
            w59=> c0_n84_w59, 
            w60=> c0_n84_w60, 
            w61=> c0_n84_w61, 
            w62=> c0_n84_w62, 
            w63=> c0_n84_w63, 
            w64=> c0_n84_w64, 
            w65=> c0_n84_w65, 
            w66=> c0_n84_w66, 
            w67=> c0_n84_w67, 
            w68=> c0_n84_w68, 
            w69=> c0_n84_w69, 
            w70=> c0_n84_w70, 
            w71=> c0_n84_w71, 
            w72=> c0_n84_w72, 
            w73=> c0_n84_w73, 
            w74=> c0_n84_w74, 
            w75=> c0_n84_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n84_y
   );           
            
neuron_inst_85: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n85_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n85_w1, 
            w2=> c0_n85_w2, 
            w3=> c0_n85_w3, 
            w4=> c0_n85_w4, 
            w5=> c0_n85_w5, 
            w6=> c0_n85_w6, 
            w7=> c0_n85_w7, 
            w8=> c0_n85_w8, 
            w9=> c0_n85_w9, 
            w10=> c0_n85_w10, 
            w11=> c0_n85_w11, 
            w12=> c0_n85_w12, 
            w13=> c0_n85_w13, 
            w14=> c0_n85_w14, 
            w15=> c0_n85_w15, 
            w16=> c0_n85_w16, 
            w17=> c0_n85_w17, 
            w18=> c0_n85_w18, 
            w19=> c0_n85_w19, 
            w20=> c0_n85_w20, 
            w21=> c0_n85_w21, 
            w22=> c0_n85_w22, 
            w23=> c0_n85_w23, 
            w24=> c0_n85_w24, 
            w25=> c0_n85_w25, 
            w26=> c0_n85_w26, 
            w27=> c0_n85_w27, 
            w28=> c0_n85_w28, 
            w29=> c0_n85_w29, 
            w30=> c0_n85_w30, 
            w31=> c0_n85_w31, 
            w32=> c0_n85_w32, 
            w33=> c0_n85_w33, 
            w34=> c0_n85_w34, 
            w35=> c0_n85_w35, 
            w36=> c0_n85_w36, 
            w37=> c0_n85_w37, 
            w38=> c0_n85_w38, 
            w39=> c0_n85_w39, 
            w40=> c0_n85_w40, 
            w41=> c0_n85_w41, 
            w42=> c0_n85_w42, 
            w43=> c0_n85_w43, 
            w44=> c0_n85_w44, 
            w45=> c0_n85_w45, 
            w46=> c0_n85_w46, 
            w47=> c0_n85_w47, 
            w48=> c0_n85_w48, 
            w49=> c0_n85_w49, 
            w50=> c0_n85_w50, 
            w51=> c0_n85_w51, 
            w52=> c0_n85_w52, 
            w53=> c0_n85_w53, 
            w54=> c0_n85_w54, 
            w55=> c0_n85_w55, 
            w56=> c0_n85_w56, 
            w57=> c0_n85_w57, 
            w58=> c0_n85_w58, 
            w59=> c0_n85_w59, 
            w60=> c0_n85_w60, 
            w61=> c0_n85_w61, 
            w62=> c0_n85_w62, 
            w63=> c0_n85_w63, 
            w64=> c0_n85_w64, 
            w65=> c0_n85_w65, 
            w66=> c0_n85_w66, 
            w67=> c0_n85_w67, 
            w68=> c0_n85_w68, 
            w69=> c0_n85_w69, 
            w70=> c0_n85_w70, 
            w71=> c0_n85_w71, 
            w72=> c0_n85_w72, 
            w73=> c0_n85_w73, 
            w74=> c0_n85_w74, 
            w75=> c0_n85_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n85_y
   );           
            
neuron_inst_86: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n86_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n86_w1, 
            w2=> c0_n86_w2, 
            w3=> c0_n86_w3, 
            w4=> c0_n86_w4, 
            w5=> c0_n86_w5, 
            w6=> c0_n86_w6, 
            w7=> c0_n86_w7, 
            w8=> c0_n86_w8, 
            w9=> c0_n86_w9, 
            w10=> c0_n86_w10, 
            w11=> c0_n86_w11, 
            w12=> c0_n86_w12, 
            w13=> c0_n86_w13, 
            w14=> c0_n86_w14, 
            w15=> c0_n86_w15, 
            w16=> c0_n86_w16, 
            w17=> c0_n86_w17, 
            w18=> c0_n86_w18, 
            w19=> c0_n86_w19, 
            w20=> c0_n86_w20, 
            w21=> c0_n86_w21, 
            w22=> c0_n86_w22, 
            w23=> c0_n86_w23, 
            w24=> c0_n86_w24, 
            w25=> c0_n86_w25, 
            w26=> c0_n86_w26, 
            w27=> c0_n86_w27, 
            w28=> c0_n86_w28, 
            w29=> c0_n86_w29, 
            w30=> c0_n86_w30, 
            w31=> c0_n86_w31, 
            w32=> c0_n86_w32, 
            w33=> c0_n86_w33, 
            w34=> c0_n86_w34, 
            w35=> c0_n86_w35, 
            w36=> c0_n86_w36, 
            w37=> c0_n86_w37, 
            w38=> c0_n86_w38, 
            w39=> c0_n86_w39, 
            w40=> c0_n86_w40, 
            w41=> c0_n86_w41, 
            w42=> c0_n86_w42, 
            w43=> c0_n86_w43, 
            w44=> c0_n86_w44, 
            w45=> c0_n86_w45, 
            w46=> c0_n86_w46, 
            w47=> c0_n86_w47, 
            w48=> c0_n86_w48, 
            w49=> c0_n86_w49, 
            w50=> c0_n86_w50, 
            w51=> c0_n86_w51, 
            w52=> c0_n86_w52, 
            w53=> c0_n86_w53, 
            w54=> c0_n86_w54, 
            w55=> c0_n86_w55, 
            w56=> c0_n86_w56, 
            w57=> c0_n86_w57, 
            w58=> c0_n86_w58, 
            w59=> c0_n86_w59, 
            w60=> c0_n86_w60, 
            w61=> c0_n86_w61, 
            w62=> c0_n86_w62, 
            w63=> c0_n86_w63, 
            w64=> c0_n86_w64, 
            w65=> c0_n86_w65, 
            w66=> c0_n86_w66, 
            w67=> c0_n86_w67, 
            w68=> c0_n86_w68, 
            w69=> c0_n86_w69, 
            w70=> c0_n86_w70, 
            w71=> c0_n86_w71, 
            w72=> c0_n86_w72, 
            w73=> c0_n86_w73, 
            w74=> c0_n86_w74, 
            w75=> c0_n86_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n86_y
   );           
            
neuron_inst_87: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n87_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n87_w1, 
            w2=> c0_n87_w2, 
            w3=> c0_n87_w3, 
            w4=> c0_n87_w4, 
            w5=> c0_n87_w5, 
            w6=> c0_n87_w6, 
            w7=> c0_n87_w7, 
            w8=> c0_n87_w8, 
            w9=> c0_n87_w9, 
            w10=> c0_n87_w10, 
            w11=> c0_n87_w11, 
            w12=> c0_n87_w12, 
            w13=> c0_n87_w13, 
            w14=> c0_n87_w14, 
            w15=> c0_n87_w15, 
            w16=> c0_n87_w16, 
            w17=> c0_n87_w17, 
            w18=> c0_n87_w18, 
            w19=> c0_n87_w19, 
            w20=> c0_n87_w20, 
            w21=> c0_n87_w21, 
            w22=> c0_n87_w22, 
            w23=> c0_n87_w23, 
            w24=> c0_n87_w24, 
            w25=> c0_n87_w25, 
            w26=> c0_n87_w26, 
            w27=> c0_n87_w27, 
            w28=> c0_n87_w28, 
            w29=> c0_n87_w29, 
            w30=> c0_n87_w30, 
            w31=> c0_n87_w31, 
            w32=> c0_n87_w32, 
            w33=> c0_n87_w33, 
            w34=> c0_n87_w34, 
            w35=> c0_n87_w35, 
            w36=> c0_n87_w36, 
            w37=> c0_n87_w37, 
            w38=> c0_n87_w38, 
            w39=> c0_n87_w39, 
            w40=> c0_n87_w40, 
            w41=> c0_n87_w41, 
            w42=> c0_n87_w42, 
            w43=> c0_n87_w43, 
            w44=> c0_n87_w44, 
            w45=> c0_n87_w45, 
            w46=> c0_n87_w46, 
            w47=> c0_n87_w47, 
            w48=> c0_n87_w48, 
            w49=> c0_n87_w49, 
            w50=> c0_n87_w50, 
            w51=> c0_n87_w51, 
            w52=> c0_n87_w52, 
            w53=> c0_n87_w53, 
            w54=> c0_n87_w54, 
            w55=> c0_n87_w55, 
            w56=> c0_n87_w56, 
            w57=> c0_n87_w57, 
            w58=> c0_n87_w58, 
            w59=> c0_n87_w59, 
            w60=> c0_n87_w60, 
            w61=> c0_n87_w61, 
            w62=> c0_n87_w62, 
            w63=> c0_n87_w63, 
            w64=> c0_n87_w64, 
            w65=> c0_n87_w65, 
            w66=> c0_n87_w66, 
            w67=> c0_n87_w67, 
            w68=> c0_n87_w68, 
            w69=> c0_n87_w69, 
            w70=> c0_n87_w70, 
            w71=> c0_n87_w71, 
            w72=> c0_n87_w72, 
            w73=> c0_n87_w73, 
            w74=> c0_n87_w74, 
            w75=> c0_n87_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n87_y
   );           
            
neuron_inst_88: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n88_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n88_w1, 
            w2=> c0_n88_w2, 
            w3=> c0_n88_w3, 
            w4=> c0_n88_w4, 
            w5=> c0_n88_w5, 
            w6=> c0_n88_w6, 
            w7=> c0_n88_w7, 
            w8=> c0_n88_w8, 
            w9=> c0_n88_w9, 
            w10=> c0_n88_w10, 
            w11=> c0_n88_w11, 
            w12=> c0_n88_w12, 
            w13=> c0_n88_w13, 
            w14=> c0_n88_w14, 
            w15=> c0_n88_w15, 
            w16=> c0_n88_w16, 
            w17=> c0_n88_w17, 
            w18=> c0_n88_w18, 
            w19=> c0_n88_w19, 
            w20=> c0_n88_w20, 
            w21=> c0_n88_w21, 
            w22=> c0_n88_w22, 
            w23=> c0_n88_w23, 
            w24=> c0_n88_w24, 
            w25=> c0_n88_w25, 
            w26=> c0_n88_w26, 
            w27=> c0_n88_w27, 
            w28=> c0_n88_w28, 
            w29=> c0_n88_w29, 
            w30=> c0_n88_w30, 
            w31=> c0_n88_w31, 
            w32=> c0_n88_w32, 
            w33=> c0_n88_w33, 
            w34=> c0_n88_w34, 
            w35=> c0_n88_w35, 
            w36=> c0_n88_w36, 
            w37=> c0_n88_w37, 
            w38=> c0_n88_w38, 
            w39=> c0_n88_w39, 
            w40=> c0_n88_w40, 
            w41=> c0_n88_w41, 
            w42=> c0_n88_w42, 
            w43=> c0_n88_w43, 
            w44=> c0_n88_w44, 
            w45=> c0_n88_w45, 
            w46=> c0_n88_w46, 
            w47=> c0_n88_w47, 
            w48=> c0_n88_w48, 
            w49=> c0_n88_w49, 
            w50=> c0_n88_w50, 
            w51=> c0_n88_w51, 
            w52=> c0_n88_w52, 
            w53=> c0_n88_w53, 
            w54=> c0_n88_w54, 
            w55=> c0_n88_w55, 
            w56=> c0_n88_w56, 
            w57=> c0_n88_w57, 
            w58=> c0_n88_w58, 
            w59=> c0_n88_w59, 
            w60=> c0_n88_w60, 
            w61=> c0_n88_w61, 
            w62=> c0_n88_w62, 
            w63=> c0_n88_w63, 
            w64=> c0_n88_w64, 
            w65=> c0_n88_w65, 
            w66=> c0_n88_w66, 
            w67=> c0_n88_w67, 
            w68=> c0_n88_w68, 
            w69=> c0_n88_w69, 
            w70=> c0_n88_w70, 
            w71=> c0_n88_w71, 
            w72=> c0_n88_w72, 
            w73=> c0_n88_w73, 
            w74=> c0_n88_w74, 
            w75=> c0_n88_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n88_y
   );           
            
neuron_inst_89: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n89_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n89_w1, 
            w2=> c0_n89_w2, 
            w3=> c0_n89_w3, 
            w4=> c0_n89_w4, 
            w5=> c0_n89_w5, 
            w6=> c0_n89_w6, 
            w7=> c0_n89_w7, 
            w8=> c0_n89_w8, 
            w9=> c0_n89_w9, 
            w10=> c0_n89_w10, 
            w11=> c0_n89_w11, 
            w12=> c0_n89_w12, 
            w13=> c0_n89_w13, 
            w14=> c0_n89_w14, 
            w15=> c0_n89_w15, 
            w16=> c0_n89_w16, 
            w17=> c0_n89_w17, 
            w18=> c0_n89_w18, 
            w19=> c0_n89_w19, 
            w20=> c0_n89_w20, 
            w21=> c0_n89_w21, 
            w22=> c0_n89_w22, 
            w23=> c0_n89_w23, 
            w24=> c0_n89_w24, 
            w25=> c0_n89_w25, 
            w26=> c0_n89_w26, 
            w27=> c0_n89_w27, 
            w28=> c0_n89_w28, 
            w29=> c0_n89_w29, 
            w30=> c0_n89_w30, 
            w31=> c0_n89_w31, 
            w32=> c0_n89_w32, 
            w33=> c0_n89_w33, 
            w34=> c0_n89_w34, 
            w35=> c0_n89_w35, 
            w36=> c0_n89_w36, 
            w37=> c0_n89_w37, 
            w38=> c0_n89_w38, 
            w39=> c0_n89_w39, 
            w40=> c0_n89_w40, 
            w41=> c0_n89_w41, 
            w42=> c0_n89_w42, 
            w43=> c0_n89_w43, 
            w44=> c0_n89_w44, 
            w45=> c0_n89_w45, 
            w46=> c0_n89_w46, 
            w47=> c0_n89_w47, 
            w48=> c0_n89_w48, 
            w49=> c0_n89_w49, 
            w50=> c0_n89_w50, 
            w51=> c0_n89_w51, 
            w52=> c0_n89_w52, 
            w53=> c0_n89_w53, 
            w54=> c0_n89_w54, 
            w55=> c0_n89_w55, 
            w56=> c0_n89_w56, 
            w57=> c0_n89_w57, 
            w58=> c0_n89_w58, 
            w59=> c0_n89_w59, 
            w60=> c0_n89_w60, 
            w61=> c0_n89_w61, 
            w62=> c0_n89_w62, 
            w63=> c0_n89_w63, 
            w64=> c0_n89_w64, 
            w65=> c0_n89_w65, 
            w66=> c0_n89_w66, 
            w67=> c0_n89_w67, 
            w68=> c0_n89_w68, 
            w69=> c0_n89_w69, 
            w70=> c0_n89_w70, 
            w71=> c0_n89_w71, 
            w72=> c0_n89_w72, 
            w73=> c0_n89_w73, 
            w74=> c0_n89_w74, 
            w75=> c0_n89_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n89_y
   );           
            
neuron_inst_90: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n90_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n90_w1, 
            w2=> c0_n90_w2, 
            w3=> c0_n90_w3, 
            w4=> c0_n90_w4, 
            w5=> c0_n90_w5, 
            w6=> c0_n90_w6, 
            w7=> c0_n90_w7, 
            w8=> c0_n90_w8, 
            w9=> c0_n90_w9, 
            w10=> c0_n90_w10, 
            w11=> c0_n90_w11, 
            w12=> c0_n90_w12, 
            w13=> c0_n90_w13, 
            w14=> c0_n90_w14, 
            w15=> c0_n90_w15, 
            w16=> c0_n90_w16, 
            w17=> c0_n90_w17, 
            w18=> c0_n90_w18, 
            w19=> c0_n90_w19, 
            w20=> c0_n90_w20, 
            w21=> c0_n90_w21, 
            w22=> c0_n90_w22, 
            w23=> c0_n90_w23, 
            w24=> c0_n90_w24, 
            w25=> c0_n90_w25, 
            w26=> c0_n90_w26, 
            w27=> c0_n90_w27, 
            w28=> c0_n90_w28, 
            w29=> c0_n90_w29, 
            w30=> c0_n90_w30, 
            w31=> c0_n90_w31, 
            w32=> c0_n90_w32, 
            w33=> c0_n90_w33, 
            w34=> c0_n90_w34, 
            w35=> c0_n90_w35, 
            w36=> c0_n90_w36, 
            w37=> c0_n90_w37, 
            w38=> c0_n90_w38, 
            w39=> c0_n90_w39, 
            w40=> c0_n90_w40, 
            w41=> c0_n90_w41, 
            w42=> c0_n90_w42, 
            w43=> c0_n90_w43, 
            w44=> c0_n90_w44, 
            w45=> c0_n90_w45, 
            w46=> c0_n90_w46, 
            w47=> c0_n90_w47, 
            w48=> c0_n90_w48, 
            w49=> c0_n90_w49, 
            w50=> c0_n90_w50, 
            w51=> c0_n90_w51, 
            w52=> c0_n90_w52, 
            w53=> c0_n90_w53, 
            w54=> c0_n90_w54, 
            w55=> c0_n90_w55, 
            w56=> c0_n90_w56, 
            w57=> c0_n90_w57, 
            w58=> c0_n90_w58, 
            w59=> c0_n90_w59, 
            w60=> c0_n90_w60, 
            w61=> c0_n90_w61, 
            w62=> c0_n90_w62, 
            w63=> c0_n90_w63, 
            w64=> c0_n90_w64, 
            w65=> c0_n90_w65, 
            w66=> c0_n90_w66, 
            w67=> c0_n90_w67, 
            w68=> c0_n90_w68, 
            w69=> c0_n90_w69, 
            w70=> c0_n90_w70, 
            w71=> c0_n90_w71, 
            w72=> c0_n90_w72, 
            w73=> c0_n90_w73, 
            w74=> c0_n90_w74, 
            w75=> c0_n90_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n90_y
   );           
            
neuron_inst_91: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n91_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n91_w1, 
            w2=> c0_n91_w2, 
            w3=> c0_n91_w3, 
            w4=> c0_n91_w4, 
            w5=> c0_n91_w5, 
            w6=> c0_n91_w6, 
            w7=> c0_n91_w7, 
            w8=> c0_n91_w8, 
            w9=> c0_n91_w9, 
            w10=> c0_n91_w10, 
            w11=> c0_n91_w11, 
            w12=> c0_n91_w12, 
            w13=> c0_n91_w13, 
            w14=> c0_n91_w14, 
            w15=> c0_n91_w15, 
            w16=> c0_n91_w16, 
            w17=> c0_n91_w17, 
            w18=> c0_n91_w18, 
            w19=> c0_n91_w19, 
            w20=> c0_n91_w20, 
            w21=> c0_n91_w21, 
            w22=> c0_n91_w22, 
            w23=> c0_n91_w23, 
            w24=> c0_n91_w24, 
            w25=> c0_n91_w25, 
            w26=> c0_n91_w26, 
            w27=> c0_n91_w27, 
            w28=> c0_n91_w28, 
            w29=> c0_n91_w29, 
            w30=> c0_n91_w30, 
            w31=> c0_n91_w31, 
            w32=> c0_n91_w32, 
            w33=> c0_n91_w33, 
            w34=> c0_n91_w34, 
            w35=> c0_n91_w35, 
            w36=> c0_n91_w36, 
            w37=> c0_n91_w37, 
            w38=> c0_n91_w38, 
            w39=> c0_n91_w39, 
            w40=> c0_n91_w40, 
            w41=> c0_n91_w41, 
            w42=> c0_n91_w42, 
            w43=> c0_n91_w43, 
            w44=> c0_n91_w44, 
            w45=> c0_n91_w45, 
            w46=> c0_n91_w46, 
            w47=> c0_n91_w47, 
            w48=> c0_n91_w48, 
            w49=> c0_n91_w49, 
            w50=> c0_n91_w50, 
            w51=> c0_n91_w51, 
            w52=> c0_n91_w52, 
            w53=> c0_n91_w53, 
            w54=> c0_n91_w54, 
            w55=> c0_n91_w55, 
            w56=> c0_n91_w56, 
            w57=> c0_n91_w57, 
            w58=> c0_n91_w58, 
            w59=> c0_n91_w59, 
            w60=> c0_n91_w60, 
            w61=> c0_n91_w61, 
            w62=> c0_n91_w62, 
            w63=> c0_n91_w63, 
            w64=> c0_n91_w64, 
            w65=> c0_n91_w65, 
            w66=> c0_n91_w66, 
            w67=> c0_n91_w67, 
            w68=> c0_n91_w68, 
            w69=> c0_n91_w69, 
            w70=> c0_n91_w70, 
            w71=> c0_n91_w71, 
            w72=> c0_n91_w72, 
            w73=> c0_n91_w73, 
            w74=> c0_n91_w74, 
            w75=> c0_n91_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n91_y
   );           
            
neuron_inst_92: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n92_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n92_w1, 
            w2=> c0_n92_w2, 
            w3=> c0_n92_w3, 
            w4=> c0_n92_w4, 
            w5=> c0_n92_w5, 
            w6=> c0_n92_w6, 
            w7=> c0_n92_w7, 
            w8=> c0_n92_w8, 
            w9=> c0_n92_w9, 
            w10=> c0_n92_w10, 
            w11=> c0_n92_w11, 
            w12=> c0_n92_w12, 
            w13=> c0_n92_w13, 
            w14=> c0_n92_w14, 
            w15=> c0_n92_w15, 
            w16=> c0_n92_w16, 
            w17=> c0_n92_w17, 
            w18=> c0_n92_w18, 
            w19=> c0_n92_w19, 
            w20=> c0_n92_w20, 
            w21=> c0_n92_w21, 
            w22=> c0_n92_w22, 
            w23=> c0_n92_w23, 
            w24=> c0_n92_w24, 
            w25=> c0_n92_w25, 
            w26=> c0_n92_w26, 
            w27=> c0_n92_w27, 
            w28=> c0_n92_w28, 
            w29=> c0_n92_w29, 
            w30=> c0_n92_w30, 
            w31=> c0_n92_w31, 
            w32=> c0_n92_w32, 
            w33=> c0_n92_w33, 
            w34=> c0_n92_w34, 
            w35=> c0_n92_w35, 
            w36=> c0_n92_w36, 
            w37=> c0_n92_w37, 
            w38=> c0_n92_w38, 
            w39=> c0_n92_w39, 
            w40=> c0_n92_w40, 
            w41=> c0_n92_w41, 
            w42=> c0_n92_w42, 
            w43=> c0_n92_w43, 
            w44=> c0_n92_w44, 
            w45=> c0_n92_w45, 
            w46=> c0_n92_w46, 
            w47=> c0_n92_w47, 
            w48=> c0_n92_w48, 
            w49=> c0_n92_w49, 
            w50=> c0_n92_w50, 
            w51=> c0_n92_w51, 
            w52=> c0_n92_w52, 
            w53=> c0_n92_w53, 
            w54=> c0_n92_w54, 
            w55=> c0_n92_w55, 
            w56=> c0_n92_w56, 
            w57=> c0_n92_w57, 
            w58=> c0_n92_w58, 
            w59=> c0_n92_w59, 
            w60=> c0_n92_w60, 
            w61=> c0_n92_w61, 
            w62=> c0_n92_w62, 
            w63=> c0_n92_w63, 
            w64=> c0_n92_w64, 
            w65=> c0_n92_w65, 
            w66=> c0_n92_w66, 
            w67=> c0_n92_w67, 
            w68=> c0_n92_w68, 
            w69=> c0_n92_w69, 
            w70=> c0_n92_w70, 
            w71=> c0_n92_w71, 
            w72=> c0_n92_w72, 
            w73=> c0_n92_w73, 
            w74=> c0_n92_w74, 
            w75=> c0_n92_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n92_y
   );           
            
neuron_inst_93: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n93_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n93_w1, 
            w2=> c0_n93_w2, 
            w3=> c0_n93_w3, 
            w4=> c0_n93_w4, 
            w5=> c0_n93_w5, 
            w6=> c0_n93_w6, 
            w7=> c0_n93_w7, 
            w8=> c0_n93_w8, 
            w9=> c0_n93_w9, 
            w10=> c0_n93_w10, 
            w11=> c0_n93_w11, 
            w12=> c0_n93_w12, 
            w13=> c0_n93_w13, 
            w14=> c0_n93_w14, 
            w15=> c0_n93_w15, 
            w16=> c0_n93_w16, 
            w17=> c0_n93_w17, 
            w18=> c0_n93_w18, 
            w19=> c0_n93_w19, 
            w20=> c0_n93_w20, 
            w21=> c0_n93_w21, 
            w22=> c0_n93_w22, 
            w23=> c0_n93_w23, 
            w24=> c0_n93_w24, 
            w25=> c0_n93_w25, 
            w26=> c0_n93_w26, 
            w27=> c0_n93_w27, 
            w28=> c0_n93_w28, 
            w29=> c0_n93_w29, 
            w30=> c0_n93_w30, 
            w31=> c0_n93_w31, 
            w32=> c0_n93_w32, 
            w33=> c0_n93_w33, 
            w34=> c0_n93_w34, 
            w35=> c0_n93_w35, 
            w36=> c0_n93_w36, 
            w37=> c0_n93_w37, 
            w38=> c0_n93_w38, 
            w39=> c0_n93_w39, 
            w40=> c0_n93_w40, 
            w41=> c0_n93_w41, 
            w42=> c0_n93_w42, 
            w43=> c0_n93_w43, 
            w44=> c0_n93_w44, 
            w45=> c0_n93_w45, 
            w46=> c0_n93_w46, 
            w47=> c0_n93_w47, 
            w48=> c0_n93_w48, 
            w49=> c0_n93_w49, 
            w50=> c0_n93_w50, 
            w51=> c0_n93_w51, 
            w52=> c0_n93_w52, 
            w53=> c0_n93_w53, 
            w54=> c0_n93_w54, 
            w55=> c0_n93_w55, 
            w56=> c0_n93_w56, 
            w57=> c0_n93_w57, 
            w58=> c0_n93_w58, 
            w59=> c0_n93_w59, 
            w60=> c0_n93_w60, 
            w61=> c0_n93_w61, 
            w62=> c0_n93_w62, 
            w63=> c0_n93_w63, 
            w64=> c0_n93_w64, 
            w65=> c0_n93_w65, 
            w66=> c0_n93_w66, 
            w67=> c0_n93_w67, 
            w68=> c0_n93_w68, 
            w69=> c0_n93_w69, 
            w70=> c0_n93_w70, 
            w71=> c0_n93_w71, 
            w72=> c0_n93_w72, 
            w73=> c0_n93_w73, 
            w74=> c0_n93_w74, 
            w75=> c0_n93_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n93_y
   );           
            
neuron_inst_94: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n94_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n94_w1, 
            w2=> c0_n94_w2, 
            w3=> c0_n94_w3, 
            w4=> c0_n94_w4, 
            w5=> c0_n94_w5, 
            w6=> c0_n94_w6, 
            w7=> c0_n94_w7, 
            w8=> c0_n94_w8, 
            w9=> c0_n94_w9, 
            w10=> c0_n94_w10, 
            w11=> c0_n94_w11, 
            w12=> c0_n94_w12, 
            w13=> c0_n94_w13, 
            w14=> c0_n94_w14, 
            w15=> c0_n94_w15, 
            w16=> c0_n94_w16, 
            w17=> c0_n94_w17, 
            w18=> c0_n94_w18, 
            w19=> c0_n94_w19, 
            w20=> c0_n94_w20, 
            w21=> c0_n94_w21, 
            w22=> c0_n94_w22, 
            w23=> c0_n94_w23, 
            w24=> c0_n94_w24, 
            w25=> c0_n94_w25, 
            w26=> c0_n94_w26, 
            w27=> c0_n94_w27, 
            w28=> c0_n94_w28, 
            w29=> c0_n94_w29, 
            w30=> c0_n94_w30, 
            w31=> c0_n94_w31, 
            w32=> c0_n94_w32, 
            w33=> c0_n94_w33, 
            w34=> c0_n94_w34, 
            w35=> c0_n94_w35, 
            w36=> c0_n94_w36, 
            w37=> c0_n94_w37, 
            w38=> c0_n94_w38, 
            w39=> c0_n94_w39, 
            w40=> c0_n94_w40, 
            w41=> c0_n94_w41, 
            w42=> c0_n94_w42, 
            w43=> c0_n94_w43, 
            w44=> c0_n94_w44, 
            w45=> c0_n94_w45, 
            w46=> c0_n94_w46, 
            w47=> c0_n94_w47, 
            w48=> c0_n94_w48, 
            w49=> c0_n94_w49, 
            w50=> c0_n94_w50, 
            w51=> c0_n94_w51, 
            w52=> c0_n94_w52, 
            w53=> c0_n94_w53, 
            w54=> c0_n94_w54, 
            w55=> c0_n94_w55, 
            w56=> c0_n94_w56, 
            w57=> c0_n94_w57, 
            w58=> c0_n94_w58, 
            w59=> c0_n94_w59, 
            w60=> c0_n94_w60, 
            w61=> c0_n94_w61, 
            w62=> c0_n94_w62, 
            w63=> c0_n94_w63, 
            w64=> c0_n94_w64, 
            w65=> c0_n94_w65, 
            w66=> c0_n94_w66, 
            w67=> c0_n94_w67, 
            w68=> c0_n94_w68, 
            w69=> c0_n94_w69, 
            w70=> c0_n94_w70, 
            w71=> c0_n94_w71, 
            w72=> c0_n94_w72, 
            w73=> c0_n94_w73, 
            w74=> c0_n94_w74, 
            w75=> c0_n94_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n94_y
   );           
            
neuron_inst_95: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n95_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n95_w1, 
            w2=> c0_n95_w2, 
            w3=> c0_n95_w3, 
            w4=> c0_n95_w4, 
            w5=> c0_n95_w5, 
            w6=> c0_n95_w6, 
            w7=> c0_n95_w7, 
            w8=> c0_n95_w8, 
            w9=> c0_n95_w9, 
            w10=> c0_n95_w10, 
            w11=> c0_n95_w11, 
            w12=> c0_n95_w12, 
            w13=> c0_n95_w13, 
            w14=> c0_n95_w14, 
            w15=> c0_n95_w15, 
            w16=> c0_n95_w16, 
            w17=> c0_n95_w17, 
            w18=> c0_n95_w18, 
            w19=> c0_n95_w19, 
            w20=> c0_n95_w20, 
            w21=> c0_n95_w21, 
            w22=> c0_n95_w22, 
            w23=> c0_n95_w23, 
            w24=> c0_n95_w24, 
            w25=> c0_n95_w25, 
            w26=> c0_n95_w26, 
            w27=> c0_n95_w27, 
            w28=> c0_n95_w28, 
            w29=> c0_n95_w29, 
            w30=> c0_n95_w30, 
            w31=> c0_n95_w31, 
            w32=> c0_n95_w32, 
            w33=> c0_n95_w33, 
            w34=> c0_n95_w34, 
            w35=> c0_n95_w35, 
            w36=> c0_n95_w36, 
            w37=> c0_n95_w37, 
            w38=> c0_n95_w38, 
            w39=> c0_n95_w39, 
            w40=> c0_n95_w40, 
            w41=> c0_n95_w41, 
            w42=> c0_n95_w42, 
            w43=> c0_n95_w43, 
            w44=> c0_n95_w44, 
            w45=> c0_n95_w45, 
            w46=> c0_n95_w46, 
            w47=> c0_n95_w47, 
            w48=> c0_n95_w48, 
            w49=> c0_n95_w49, 
            w50=> c0_n95_w50, 
            w51=> c0_n95_w51, 
            w52=> c0_n95_w52, 
            w53=> c0_n95_w53, 
            w54=> c0_n95_w54, 
            w55=> c0_n95_w55, 
            w56=> c0_n95_w56, 
            w57=> c0_n95_w57, 
            w58=> c0_n95_w58, 
            w59=> c0_n95_w59, 
            w60=> c0_n95_w60, 
            w61=> c0_n95_w61, 
            w62=> c0_n95_w62, 
            w63=> c0_n95_w63, 
            w64=> c0_n95_w64, 
            w65=> c0_n95_w65, 
            w66=> c0_n95_w66, 
            w67=> c0_n95_w67, 
            w68=> c0_n95_w68, 
            w69=> c0_n95_w69, 
            w70=> c0_n95_w70, 
            w71=> c0_n95_w71, 
            w72=> c0_n95_w72, 
            w73=> c0_n95_w73, 
            w74=> c0_n95_w74, 
            w75=> c0_n95_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n95_y
   );           
            
neuron_inst_96: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n96_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n96_w1, 
            w2=> c0_n96_w2, 
            w3=> c0_n96_w3, 
            w4=> c0_n96_w4, 
            w5=> c0_n96_w5, 
            w6=> c0_n96_w6, 
            w7=> c0_n96_w7, 
            w8=> c0_n96_w8, 
            w9=> c0_n96_w9, 
            w10=> c0_n96_w10, 
            w11=> c0_n96_w11, 
            w12=> c0_n96_w12, 
            w13=> c0_n96_w13, 
            w14=> c0_n96_w14, 
            w15=> c0_n96_w15, 
            w16=> c0_n96_w16, 
            w17=> c0_n96_w17, 
            w18=> c0_n96_w18, 
            w19=> c0_n96_w19, 
            w20=> c0_n96_w20, 
            w21=> c0_n96_w21, 
            w22=> c0_n96_w22, 
            w23=> c0_n96_w23, 
            w24=> c0_n96_w24, 
            w25=> c0_n96_w25, 
            w26=> c0_n96_w26, 
            w27=> c0_n96_w27, 
            w28=> c0_n96_w28, 
            w29=> c0_n96_w29, 
            w30=> c0_n96_w30, 
            w31=> c0_n96_w31, 
            w32=> c0_n96_w32, 
            w33=> c0_n96_w33, 
            w34=> c0_n96_w34, 
            w35=> c0_n96_w35, 
            w36=> c0_n96_w36, 
            w37=> c0_n96_w37, 
            w38=> c0_n96_w38, 
            w39=> c0_n96_w39, 
            w40=> c0_n96_w40, 
            w41=> c0_n96_w41, 
            w42=> c0_n96_w42, 
            w43=> c0_n96_w43, 
            w44=> c0_n96_w44, 
            w45=> c0_n96_w45, 
            w46=> c0_n96_w46, 
            w47=> c0_n96_w47, 
            w48=> c0_n96_w48, 
            w49=> c0_n96_w49, 
            w50=> c0_n96_w50, 
            w51=> c0_n96_w51, 
            w52=> c0_n96_w52, 
            w53=> c0_n96_w53, 
            w54=> c0_n96_w54, 
            w55=> c0_n96_w55, 
            w56=> c0_n96_w56, 
            w57=> c0_n96_w57, 
            w58=> c0_n96_w58, 
            w59=> c0_n96_w59, 
            w60=> c0_n96_w60, 
            w61=> c0_n96_w61, 
            w62=> c0_n96_w62, 
            w63=> c0_n96_w63, 
            w64=> c0_n96_w64, 
            w65=> c0_n96_w65, 
            w66=> c0_n96_w66, 
            w67=> c0_n96_w67, 
            w68=> c0_n96_w68, 
            w69=> c0_n96_w69, 
            w70=> c0_n96_w70, 
            w71=> c0_n96_w71, 
            w72=> c0_n96_w72, 
            w73=> c0_n96_w73, 
            w74=> c0_n96_w74, 
            w75=> c0_n96_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n96_y
   );           
            
neuron_inst_97: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n97_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n97_w1, 
            w2=> c0_n97_w2, 
            w3=> c0_n97_w3, 
            w4=> c0_n97_w4, 
            w5=> c0_n97_w5, 
            w6=> c0_n97_w6, 
            w7=> c0_n97_w7, 
            w8=> c0_n97_w8, 
            w9=> c0_n97_w9, 
            w10=> c0_n97_w10, 
            w11=> c0_n97_w11, 
            w12=> c0_n97_w12, 
            w13=> c0_n97_w13, 
            w14=> c0_n97_w14, 
            w15=> c0_n97_w15, 
            w16=> c0_n97_w16, 
            w17=> c0_n97_w17, 
            w18=> c0_n97_w18, 
            w19=> c0_n97_w19, 
            w20=> c0_n97_w20, 
            w21=> c0_n97_w21, 
            w22=> c0_n97_w22, 
            w23=> c0_n97_w23, 
            w24=> c0_n97_w24, 
            w25=> c0_n97_w25, 
            w26=> c0_n97_w26, 
            w27=> c0_n97_w27, 
            w28=> c0_n97_w28, 
            w29=> c0_n97_w29, 
            w30=> c0_n97_w30, 
            w31=> c0_n97_w31, 
            w32=> c0_n97_w32, 
            w33=> c0_n97_w33, 
            w34=> c0_n97_w34, 
            w35=> c0_n97_w35, 
            w36=> c0_n97_w36, 
            w37=> c0_n97_w37, 
            w38=> c0_n97_w38, 
            w39=> c0_n97_w39, 
            w40=> c0_n97_w40, 
            w41=> c0_n97_w41, 
            w42=> c0_n97_w42, 
            w43=> c0_n97_w43, 
            w44=> c0_n97_w44, 
            w45=> c0_n97_w45, 
            w46=> c0_n97_w46, 
            w47=> c0_n97_w47, 
            w48=> c0_n97_w48, 
            w49=> c0_n97_w49, 
            w50=> c0_n97_w50, 
            w51=> c0_n97_w51, 
            w52=> c0_n97_w52, 
            w53=> c0_n97_w53, 
            w54=> c0_n97_w54, 
            w55=> c0_n97_w55, 
            w56=> c0_n97_w56, 
            w57=> c0_n97_w57, 
            w58=> c0_n97_w58, 
            w59=> c0_n97_w59, 
            w60=> c0_n97_w60, 
            w61=> c0_n97_w61, 
            w62=> c0_n97_w62, 
            w63=> c0_n97_w63, 
            w64=> c0_n97_w64, 
            w65=> c0_n97_w65, 
            w66=> c0_n97_w66, 
            w67=> c0_n97_w67, 
            w68=> c0_n97_w68, 
            w69=> c0_n97_w69, 
            w70=> c0_n97_w70, 
            w71=> c0_n97_w71, 
            w72=> c0_n97_w72, 
            w73=> c0_n97_w73, 
            w74=> c0_n97_w74, 
            w75=> c0_n97_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n97_y
   );           
            
neuron_inst_98: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n98_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n98_w1, 
            w2=> c0_n98_w2, 
            w3=> c0_n98_w3, 
            w4=> c0_n98_w4, 
            w5=> c0_n98_w5, 
            w6=> c0_n98_w6, 
            w7=> c0_n98_w7, 
            w8=> c0_n98_w8, 
            w9=> c0_n98_w9, 
            w10=> c0_n98_w10, 
            w11=> c0_n98_w11, 
            w12=> c0_n98_w12, 
            w13=> c0_n98_w13, 
            w14=> c0_n98_w14, 
            w15=> c0_n98_w15, 
            w16=> c0_n98_w16, 
            w17=> c0_n98_w17, 
            w18=> c0_n98_w18, 
            w19=> c0_n98_w19, 
            w20=> c0_n98_w20, 
            w21=> c0_n98_w21, 
            w22=> c0_n98_w22, 
            w23=> c0_n98_w23, 
            w24=> c0_n98_w24, 
            w25=> c0_n98_w25, 
            w26=> c0_n98_w26, 
            w27=> c0_n98_w27, 
            w28=> c0_n98_w28, 
            w29=> c0_n98_w29, 
            w30=> c0_n98_w30, 
            w31=> c0_n98_w31, 
            w32=> c0_n98_w32, 
            w33=> c0_n98_w33, 
            w34=> c0_n98_w34, 
            w35=> c0_n98_w35, 
            w36=> c0_n98_w36, 
            w37=> c0_n98_w37, 
            w38=> c0_n98_w38, 
            w39=> c0_n98_w39, 
            w40=> c0_n98_w40, 
            w41=> c0_n98_w41, 
            w42=> c0_n98_w42, 
            w43=> c0_n98_w43, 
            w44=> c0_n98_w44, 
            w45=> c0_n98_w45, 
            w46=> c0_n98_w46, 
            w47=> c0_n98_w47, 
            w48=> c0_n98_w48, 
            w49=> c0_n98_w49, 
            w50=> c0_n98_w50, 
            w51=> c0_n98_w51, 
            w52=> c0_n98_w52, 
            w53=> c0_n98_w53, 
            w54=> c0_n98_w54, 
            w55=> c0_n98_w55, 
            w56=> c0_n98_w56, 
            w57=> c0_n98_w57, 
            w58=> c0_n98_w58, 
            w59=> c0_n98_w59, 
            w60=> c0_n98_w60, 
            w61=> c0_n98_w61, 
            w62=> c0_n98_w62, 
            w63=> c0_n98_w63, 
            w64=> c0_n98_w64, 
            w65=> c0_n98_w65, 
            w66=> c0_n98_w66, 
            w67=> c0_n98_w67, 
            w68=> c0_n98_w68, 
            w69=> c0_n98_w69, 
            w70=> c0_n98_w70, 
            w71=> c0_n98_w71, 
            w72=> c0_n98_w72, 
            w73=> c0_n98_w73, 
            w74=> c0_n98_w74, 
            w75=> c0_n98_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n98_y
   );           
            
neuron_inst_99: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_75n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c0_n99_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            w1=> c0_n99_w1, 
            w2=> c0_n99_w2, 
            w3=> c0_n99_w3, 
            w4=> c0_n99_w4, 
            w5=> c0_n99_w5, 
            w6=> c0_n99_w6, 
            w7=> c0_n99_w7, 
            w8=> c0_n99_w8, 
            w9=> c0_n99_w9, 
            w10=> c0_n99_w10, 
            w11=> c0_n99_w11, 
            w12=> c0_n99_w12, 
            w13=> c0_n99_w13, 
            w14=> c0_n99_w14, 
            w15=> c0_n99_w15, 
            w16=> c0_n99_w16, 
            w17=> c0_n99_w17, 
            w18=> c0_n99_w18, 
            w19=> c0_n99_w19, 
            w20=> c0_n99_w20, 
            w21=> c0_n99_w21, 
            w22=> c0_n99_w22, 
            w23=> c0_n99_w23, 
            w24=> c0_n99_w24, 
            w25=> c0_n99_w25, 
            w26=> c0_n99_w26, 
            w27=> c0_n99_w27, 
            w28=> c0_n99_w28, 
            w29=> c0_n99_w29, 
            w30=> c0_n99_w30, 
            w31=> c0_n99_w31, 
            w32=> c0_n99_w32, 
            w33=> c0_n99_w33, 
            w34=> c0_n99_w34, 
            w35=> c0_n99_w35, 
            w36=> c0_n99_w36, 
            w37=> c0_n99_w37, 
            w38=> c0_n99_w38, 
            w39=> c0_n99_w39, 
            w40=> c0_n99_w40, 
            w41=> c0_n99_w41, 
            w42=> c0_n99_w42, 
            w43=> c0_n99_w43, 
            w44=> c0_n99_w44, 
            w45=> c0_n99_w45, 
            w46=> c0_n99_w46, 
            w47=> c0_n99_w47, 
            w48=> c0_n99_w48, 
            w49=> c0_n99_w49, 
            w50=> c0_n99_w50, 
            w51=> c0_n99_w51, 
            w52=> c0_n99_w52, 
            w53=> c0_n99_w53, 
            w54=> c0_n99_w54, 
            w55=> c0_n99_w55, 
            w56=> c0_n99_w56, 
            w57=> c0_n99_w57, 
            w58=> c0_n99_w58, 
            w59=> c0_n99_w59, 
            w60=> c0_n99_w60, 
            w61=> c0_n99_w61, 
            w62=> c0_n99_w62, 
            w63=> c0_n99_w63, 
            w64=> c0_n99_w64, 
            w65=> c0_n99_w65, 
            w66=> c0_n99_w66, 
            w67=> c0_n99_w67, 
            w68=> c0_n99_w68, 
            w69=> c0_n99_w69, 
            w70=> c0_n99_w70, 
            w71=> c0_n99_w71, 
            w72=> c0_n99_w72, 
            w73=> c0_n99_w73, 
            w74=> c0_n99_w74, 
            w75=> c0_n99_w75, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c0_n99_y
   );           
             
END ARCHITECTURE;
