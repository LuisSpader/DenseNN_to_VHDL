LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY  camada1_Leaky_ReLU_30neuron_8bits_100n_signed IS
  PORT (
    clk, rst: IN STD_LOGIC;
    c1_n0_bias, c1_n1_bias, c1_n2_bias, c1_n3_bias, c1_n4_bias, c1_n5_bias, c1_n6_bias, c1_n7_bias, c1_n8_bias, c1_n9_bias, c1_n10_bias, c1_n11_bias, c1_n12_bias, c1_n13_bias, c1_n14_bias, c1_n15_bias, c1_n16_bias, c1_n17_bias, c1_n18_bias, c1_n19_bias, c1_n20_bias, c1_n21_bias, c1_n22_bias, c1_n23_bias, c1_n24_bias, c1_n25_bias, c1_n26_bias, c1_n27_bias, c1_n28_bias, c1_n29_bias, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, c1_n0_w1, c1_n0_w2, c1_n0_w3, c1_n0_w4, c1_n0_w5, c1_n0_w6, c1_n0_w7, c1_n0_w8, c1_n0_w9, c1_n0_w10, c1_n0_w11, c1_n0_w12, c1_n0_w13, c1_n0_w14, c1_n0_w15, c1_n0_w16, c1_n0_w17, c1_n0_w18, c1_n0_w19, c1_n0_w20, c1_n0_w21, c1_n0_w22, c1_n0_w23, c1_n0_w24, c1_n0_w25, c1_n0_w26, c1_n0_w27, c1_n0_w28, c1_n0_w29, c1_n0_w30, c1_n0_w31, c1_n0_w32, c1_n0_w33, c1_n0_w34, c1_n0_w35, c1_n0_w36, c1_n0_w37, c1_n0_w38, c1_n0_w39, c1_n0_w40, c1_n0_w41, c1_n0_w42, c1_n0_w43, c1_n0_w44, c1_n0_w45, c1_n0_w46, c1_n0_w47, c1_n0_w48, c1_n0_w49, c1_n0_w50, c1_n0_w51, c1_n0_w52, c1_n0_w53, c1_n0_w54, c1_n0_w55, c1_n0_w56, c1_n0_w57, c1_n0_w58, c1_n0_w59, c1_n0_w60, c1_n0_w61, c1_n0_w62, c1_n0_w63, c1_n0_w64, c1_n0_w65, c1_n0_w66, c1_n0_w67, c1_n0_w68, c1_n0_w69, c1_n0_w70, c1_n0_w71, c1_n0_w72, c1_n0_w73, c1_n0_w74, c1_n0_w75, c1_n0_w76, c1_n0_w77, c1_n0_w78, c1_n0_w79, c1_n0_w80, c1_n0_w81, c1_n0_w82, c1_n0_w83, c1_n0_w84, c1_n0_w85, c1_n0_w86, c1_n0_w87, c1_n0_w88, c1_n0_w89, c1_n0_w90, c1_n0_w91, c1_n0_w92, c1_n0_w93, c1_n0_w94, c1_n0_w95, c1_n0_w96, c1_n0_w97, c1_n0_w98, c1_n0_w99, c1_n0_w100, c1_n1_w1, c1_n1_w2, c1_n1_w3, c1_n1_w4, c1_n1_w5, c1_n1_w6, c1_n1_w7, c1_n1_w8, c1_n1_w9, c1_n1_w10, c1_n1_w11, c1_n1_w12, c1_n1_w13, c1_n1_w14, c1_n1_w15, c1_n1_w16, c1_n1_w17, c1_n1_w18, c1_n1_w19, c1_n1_w20, c1_n1_w21, c1_n1_w22, c1_n1_w23, c1_n1_w24, c1_n1_w25, c1_n1_w26, c1_n1_w27, c1_n1_w28, c1_n1_w29, c1_n1_w30, c1_n1_w31, c1_n1_w32, c1_n1_w33, c1_n1_w34, c1_n1_w35, c1_n1_w36, c1_n1_w37, c1_n1_w38, c1_n1_w39, c1_n1_w40, c1_n1_w41, c1_n1_w42, c1_n1_w43, c1_n1_w44, c1_n1_w45, c1_n1_w46, c1_n1_w47, c1_n1_w48, c1_n1_w49, c1_n1_w50, c1_n1_w51, c1_n1_w52, c1_n1_w53, c1_n1_w54, c1_n1_w55, c1_n1_w56, c1_n1_w57, c1_n1_w58, c1_n1_w59, c1_n1_w60, c1_n1_w61, c1_n1_w62, c1_n1_w63, c1_n1_w64, c1_n1_w65, c1_n1_w66, c1_n1_w67, c1_n1_w68, c1_n1_w69, c1_n1_w70, c1_n1_w71, c1_n1_w72, c1_n1_w73, c1_n1_w74, c1_n1_w75, c1_n1_w76, c1_n1_w77, c1_n1_w78, c1_n1_w79, c1_n1_w80, c1_n1_w81, c1_n1_w82, c1_n1_w83, c1_n1_w84, c1_n1_w85, c1_n1_w86, c1_n1_w87, c1_n1_w88, c1_n1_w89, c1_n1_w90, c1_n1_w91, c1_n1_w92, c1_n1_w93, c1_n1_w94, c1_n1_w95, c1_n1_w96, c1_n1_w97, c1_n1_w98, c1_n1_w99, c1_n1_w100, c1_n2_w1, c1_n2_w2, c1_n2_w3, c1_n2_w4, c1_n2_w5, c1_n2_w6, c1_n2_w7, c1_n2_w8, c1_n2_w9, c1_n2_w10, c1_n2_w11, c1_n2_w12, c1_n2_w13, c1_n2_w14, c1_n2_w15, c1_n2_w16, c1_n2_w17, c1_n2_w18, c1_n2_w19, c1_n2_w20, c1_n2_w21, c1_n2_w22, c1_n2_w23, c1_n2_w24, c1_n2_w25, c1_n2_w26, c1_n2_w27, c1_n2_w28, c1_n2_w29, c1_n2_w30, c1_n2_w31, c1_n2_w32, c1_n2_w33, c1_n2_w34, c1_n2_w35, c1_n2_w36, c1_n2_w37, c1_n2_w38, c1_n2_w39, c1_n2_w40, c1_n2_w41, c1_n2_w42, c1_n2_w43, c1_n2_w44, c1_n2_w45, c1_n2_w46, c1_n2_w47, c1_n2_w48, c1_n2_w49, c1_n2_w50, c1_n2_w51, c1_n2_w52, c1_n2_w53, c1_n2_w54, c1_n2_w55, c1_n2_w56, c1_n2_w57, c1_n2_w58, c1_n2_w59, c1_n2_w60, c1_n2_w61, c1_n2_w62, c1_n2_w63, c1_n2_w64, c1_n2_w65, c1_n2_w66, c1_n2_w67, c1_n2_w68, c1_n2_w69, c1_n2_w70, c1_n2_w71, c1_n2_w72, c1_n2_w73, c1_n2_w74, c1_n2_w75, c1_n2_w76, c1_n2_w77, c1_n2_w78, c1_n2_w79, c1_n2_w80, c1_n2_w81, c1_n2_w82, c1_n2_w83, c1_n2_w84, c1_n2_w85, c1_n2_w86, c1_n2_w87, c1_n2_w88, c1_n2_w89, c1_n2_w90, c1_n2_w91, c1_n2_w92, c1_n2_w93, c1_n2_w94, c1_n2_w95, c1_n2_w96, c1_n2_w97, c1_n2_w98, c1_n2_w99, c1_n2_w100, c1_n3_w1, c1_n3_w2, c1_n3_w3, c1_n3_w4, c1_n3_w5, c1_n3_w6, c1_n3_w7, c1_n3_w8, c1_n3_w9, c1_n3_w10, c1_n3_w11, c1_n3_w12, c1_n3_w13, c1_n3_w14, c1_n3_w15, c1_n3_w16, c1_n3_w17, c1_n3_w18, c1_n3_w19, c1_n3_w20, c1_n3_w21, c1_n3_w22, c1_n3_w23, c1_n3_w24, c1_n3_w25, c1_n3_w26, c1_n3_w27, c1_n3_w28, c1_n3_w29, c1_n3_w30, c1_n3_w31, c1_n3_w32, c1_n3_w33, c1_n3_w34, c1_n3_w35, c1_n3_w36, c1_n3_w37, c1_n3_w38, c1_n3_w39, c1_n3_w40, c1_n3_w41, c1_n3_w42, c1_n3_w43, c1_n3_w44, c1_n3_w45, c1_n3_w46, c1_n3_w47, c1_n3_w48, c1_n3_w49, c1_n3_w50, c1_n3_w51, c1_n3_w52, c1_n3_w53, c1_n3_w54, c1_n3_w55, c1_n3_w56, c1_n3_w57, c1_n3_w58, c1_n3_w59, c1_n3_w60, c1_n3_w61, c1_n3_w62, c1_n3_w63, c1_n3_w64, c1_n3_w65, c1_n3_w66, c1_n3_w67, c1_n3_w68, c1_n3_w69, c1_n3_w70, c1_n3_w71, c1_n3_w72, c1_n3_w73, c1_n3_w74, c1_n3_w75, c1_n3_w76, c1_n3_w77, c1_n3_w78, c1_n3_w79, c1_n3_w80, c1_n3_w81, c1_n3_w82, c1_n3_w83, c1_n3_w84, c1_n3_w85, c1_n3_w86, c1_n3_w87, c1_n3_w88, c1_n3_w89, c1_n3_w90, c1_n3_w91, c1_n3_w92, c1_n3_w93, c1_n3_w94, c1_n3_w95, c1_n3_w96, c1_n3_w97, c1_n3_w98, c1_n3_w99, c1_n3_w100, c1_n4_w1, c1_n4_w2, c1_n4_w3, c1_n4_w4, c1_n4_w5, c1_n4_w6, c1_n4_w7, c1_n4_w8, c1_n4_w9, c1_n4_w10, c1_n4_w11, c1_n4_w12, c1_n4_w13, c1_n4_w14, c1_n4_w15, c1_n4_w16, c1_n4_w17, c1_n4_w18, c1_n4_w19, c1_n4_w20, c1_n4_w21, c1_n4_w22, c1_n4_w23, c1_n4_w24, c1_n4_w25, c1_n4_w26, c1_n4_w27, c1_n4_w28, c1_n4_w29, c1_n4_w30, c1_n4_w31, c1_n4_w32, c1_n4_w33, c1_n4_w34, c1_n4_w35, c1_n4_w36, c1_n4_w37, c1_n4_w38, c1_n4_w39, c1_n4_w40, c1_n4_w41, c1_n4_w42, c1_n4_w43, c1_n4_w44, c1_n4_w45, c1_n4_w46, c1_n4_w47, c1_n4_w48, c1_n4_w49, c1_n4_w50, c1_n4_w51, c1_n4_w52, c1_n4_w53, c1_n4_w54, c1_n4_w55, c1_n4_w56, c1_n4_w57, c1_n4_w58, c1_n4_w59, c1_n4_w60, c1_n4_w61, c1_n4_w62, c1_n4_w63, c1_n4_w64, c1_n4_w65, c1_n4_w66, c1_n4_w67, c1_n4_w68, c1_n4_w69, c1_n4_w70, c1_n4_w71, c1_n4_w72, c1_n4_w73, c1_n4_w74, c1_n4_w75, c1_n4_w76, c1_n4_w77, c1_n4_w78, c1_n4_w79, c1_n4_w80, c1_n4_w81, c1_n4_w82, c1_n4_w83, c1_n4_w84, c1_n4_w85, c1_n4_w86, c1_n4_w87, c1_n4_w88, c1_n4_w89, c1_n4_w90, c1_n4_w91, c1_n4_w92, c1_n4_w93, c1_n4_w94, c1_n4_w95, c1_n4_w96, c1_n4_w97, c1_n4_w98, c1_n4_w99, c1_n4_w100, c1_n5_w1, c1_n5_w2, c1_n5_w3, c1_n5_w4, c1_n5_w5, c1_n5_w6, c1_n5_w7, c1_n5_w8, c1_n5_w9, c1_n5_w10, c1_n5_w11, c1_n5_w12, c1_n5_w13, c1_n5_w14, c1_n5_w15, c1_n5_w16, c1_n5_w17, c1_n5_w18, c1_n5_w19, c1_n5_w20, c1_n5_w21, c1_n5_w22, c1_n5_w23, c1_n5_w24, c1_n5_w25, c1_n5_w26, c1_n5_w27, c1_n5_w28, c1_n5_w29, c1_n5_w30, c1_n5_w31, c1_n5_w32, c1_n5_w33, c1_n5_w34, c1_n5_w35, c1_n5_w36, c1_n5_w37, c1_n5_w38, c1_n5_w39, c1_n5_w40, c1_n5_w41, c1_n5_w42, c1_n5_w43, c1_n5_w44, c1_n5_w45, c1_n5_w46, c1_n5_w47, c1_n5_w48, c1_n5_w49, c1_n5_w50, c1_n5_w51, c1_n5_w52, c1_n5_w53, c1_n5_w54, c1_n5_w55, c1_n5_w56, c1_n5_w57, c1_n5_w58, c1_n5_w59, c1_n5_w60, c1_n5_w61, c1_n5_w62, c1_n5_w63, c1_n5_w64, c1_n5_w65, c1_n5_w66, c1_n5_w67, c1_n5_w68, c1_n5_w69, c1_n5_w70, c1_n5_w71, c1_n5_w72, c1_n5_w73, c1_n5_w74, c1_n5_w75, c1_n5_w76, c1_n5_w77, c1_n5_w78, c1_n5_w79, c1_n5_w80, c1_n5_w81, c1_n5_w82, c1_n5_w83, c1_n5_w84, c1_n5_w85, c1_n5_w86, c1_n5_w87, c1_n5_w88, c1_n5_w89, c1_n5_w90, c1_n5_w91, c1_n5_w92, c1_n5_w93, c1_n5_w94, c1_n5_w95, c1_n5_w96, c1_n5_w97, c1_n5_w98, c1_n5_w99, c1_n5_w100, c1_n6_w1, c1_n6_w2, c1_n6_w3, c1_n6_w4, c1_n6_w5, c1_n6_w6, c1_n6_w7, c1_n6_w8, c1_n6_w9, c1_n6_w10, c1_n6_w11, c1_n6_w12, c1_n6_w13, c1_n6_w14, c1_n6_w15, c1_n6_w16, c1_n6_w17, c1_n6_w18, c1_n6_w19, c1_n6_w20, c1_n6_w21, c1_n6_w22, c1_n6_w23, c1_n6_w24, c1_n6_w25, c1_n6_w26, c1_n6_w27, c1_n6_w28, c1_n6_w29, c1_n6_w30, c1_n6_w31, c1_n6_w32, c1_n6_w33, c1_n6_w34, c1_n6_w35, c1_n6_w36, c1_n6_w37, c1_n6_w38, c1_n6_w39, c1_n6_w40, c1_n6_w41, c1_n6_w42, c1_n6_w43, c1_n6_w44, c1_n6_w45, c1_n6_w46, c1_n6_w47, c1_n6_w48, c1_n6_w49, c1_n6_w50, c1_n6_w51, c1_n6_w52, c1_n6_w53, c1_n6_w54, c1_n6_w55, c1_n6_w56, c1_n6_w57, c1_n6_w58, c1_n6_w59, c1_n6_w60, c1_n6_w61, c1_n6_w62, c1_n6_w63, c1_n6_w64, c1_n6_w65, c1_n6_w66, c1_n6_w67, c1_n6_w68, c1_n6_w69, c1_n6_w70, c1_n6_w71, c1_n6_w72, c1_n6_w73, c1_n6_w74, c1_n6_w75, c1_n6_w76, c1_n6_w77, c1_n6_w78, c1_n6_w79, c1_n6_w80, c1_n6_w81, c1_n6_w82, c1_n6_w83, c1_n6_w84, c1_n6_w85, c1_n6_w86, c1_n6_w87, c1_n6_w88, c1_n6_w89, c1_n6_w90, c1_n6_w91, c1_n6_w92, c1_n6_w93, c1_n6_w94, c1_n6_w95, c1_n6_w96, c1_n6_w97, c1_n6_w98, c1_n6_w99, c1_n6_w100, c1_n7_w1, c1_n7_w2, c1_n7_w3, c1_n7_w4, c1_n7_w5, c1_n7_w6, c1_n7_w7, c1_n7_w8, c1_n7_w9, c1_n7_w10, c1_n7_w11, c1_n7_w12, c1_n7_w13, c1_n7_w14, c1_n7_w15, c1_n7_w16, c1_n7_w17, c1_n7_w18, c1_n7_w19, c1_n7_w20, c1_n7_w21, c1_n7_w22, c1_n7_w23, c1_n7_w24, c1_n7_w25, c1_n7_w26, c1_n7_w27, c1_n7_w28, c1_n7_w29, c1_n7_w30, c1_n7_w31, c1_n7_w32, c1_n7_w33, c1_n7_w34, c1_n7_w35, c1_n7_w36, c1_n7_w37, c1_n7_w38, c1_n7_w39, c1_n7_w40, c1_n7_w41, c1_n7_w42, c1_n7_w43, c1_n7_w44, c1_n7_w45, c1_n7_w46, c1_n7_w47, c1_n7_w48, c1_n7_w49, c1_n7_w50, c1_n7_w51, c1_n7_w52, c1_n7_w53, c1_n7_w54, c1_n7_w55, c1_n7_w56, c1_n7_w57, c1_n7_w58, c1_n7_w59, c1_n7_w60, c1_n7_w61, c1_n7_w62, c1_n7_w63, c1_n7_w64, c1_n7_w65, c1_n7_w66, c1_n7_w67, c1_n7_w68, c1_n7_w69, c1_n7_w70, c1_n7_w71, c1_n7_w72, c1_n7_w73, c1_n7_w74, c1_n7_w75, c1_n7_w76, c1_n7_w77, c1_n7_w78, c1_n7_w79, c1_n7_w80, c1_n7_w81, c1_n7_w82, c1_n7_w83, c1_n7_w84, c1_n7_w85, c1_n7_w86, c1_n7_w87, c1_n7_w88, c1_n7_w89, c1_n7_w90, c1_n7_w91, c1_n7_w92, c1_n7_w93, c1_n7_w94, c1_n7_w95, c1_n7_w96, c1_n7_w97, c1_n7_w98, c1_n7_w99, c1_n7_w100, c1_n8_w1, c1_n8_w2, c1_n8_w3, c1_n8_w4, c1_n8_w5, c1_n8_w6, c1_n8_w7, c1_n8_w8, c1_n8_w9, c1_n8_w10, c1_n8_w11, c1_n8_w12, c1_n8_w13, c1_n8_w14, c1_n8_w15, c1_n8_w16, c1_n8_w17, c1_n8_w18, c1_n8_w19, c1_n8_w20, c1_n8_w21, c1_n8_w22, c1_n8_w23, c1_n8_w24, c1_n8_w25, c1_n8_w26, c1_n8_w27, c1_n8_w28, c1_n8_w29, c1_n8_w30, c1_n8_w31, c1_n8_w32, c1_n8_w33, c1_n8_w34, c1_n8_w35, c1_n8_w36, c1_n8_w37, c1_n8_w38, c1_n8_w39, c1_n8_w40, c1_n8_w41, c1_n8_w42, c1_n8_w43, c1_n8_w44, c1_n8_w45, c1_n8_w46, c1_n8_w47, c1_n8_w48, c1_n8_w49, c1_n8_w50, c1_n8_w51, c1_n8_w52, c1_n8_w53, c1_n8_w54, c1_n8_w55, c1_n8_w56, c1_n8_w57, c1_n8_w58, c1_n8_w59, c1_n8_w60, c1_n8_w61, c1_n8_w62, c1_n8_w63, c1_n8_w64, c1_n8_w65, c1_n8_w66, c1_n8_w67, c1_n8_w68, c1_n8_w69, c1_n8_w70, c1_n8_w71, c1_n8_w72, c1_n8_w73, c1_n8_w74, c1_n8_w75, c1_n8_w76, c1_n8_w77, c1_n8_w78, c1_n8_w79, c1_n8_w80, c1_n8_w81, c1_n8_w82, c1_n8_w83, c1_n8_w84, c1_n8_w85, c1_n8_w86, c1_n8_w87, c1_n8_w88, c1_n8_w89, c1_n8_w90, c1_n8_w91, c1_n8_w92, c1_n8_w93, c1_n8_w94, c1_n8_w95, c1_n8_w96, c1_n8_w97, c1_n8_w98, c1_n8_w99, c1_n8_w100, c1_n9_w1, c1_n9_w2, c1_n9_w3, c1_n9_w4, c1_n9_w5, c1_n9_w6, c1_n9_w7, c1_n9_w8, c1_n9_w9, c1_n9_w10, c1_n9_w11, c1_n9_w12, c1_n9_w13, c1_n9_w14, c1_n9_w15, c1_n9_w16, c1_n9_w17, c1_n9_w18, c1_n9_w19, c1_n9_w20, c1_n9_w21, c1_n9_w22, c1_n9_w23, c1_n9_w24, c1_n9_w25, c1_n9_w26, c1_n9_w27, c1_n9_w28, c1_n9_w29, c1_n9_w30, c1_n9_w31, c1_n9_w32, c1_n9_w33, c1_n9_w34, c1_n9_w35, c1_n9_w36, c1_n9_w37, c1_n9_w38, c1_n9_w39, c1_n9_w40, c1_n9_w41, c1_n9_w42, c1_n9_w43, c1_n9_w44, c1_n9_w45, c1_n9_w46, c1_n9_w47, c1_n9_w48, c1_n9_w49, c1_n9_w50, c1_n9_w51, c1_n9_w52, c1_n9_w53, c1_n9_w54, c1_n9_w55, c1_n9_w56, c1_n9_w57, c1_n9_w58, c1_n9_w59, c1_n9_w60, c1_n9_w61, c1_n9_w62, c1_n9_w63, c1_n9_w64, c1_n9_w65, c1_n9_w66, c1_n9_w67, c1_n9_w68, c1_n9_w69, c1_n9_w70, c1_n9_w71, c1_n9_w72, c1_n9_w73, c1_n9_w74, c1_n9_w75, c1_n9_w76, c1_n9_w77, c1_n9_w78, c1_n9_w79, c1_n9_w80, c1_n9_w81, c1_n9_w82, c1_n9_w83, c1_n9_w84, c1_n9_w85, c1_n9_w86, c1_n9_w87, c1_n9_w88, c1_n9_w89, c1_n9_w90, c1_n9_w91, c1_n9_w92, c1_n9_w93, c1_n9_w94, c1_n9_w95, c1_n9_w96, c1_n9_w97, c1_n9_w98, c1_n9_w99, c1_n9_w100, c1_n10_w1, c1_n10_w2, c1_n10_w3, c1_n10_w4, c1_n10_w5, c1_n10_w6, c1_n10_w7, c1_n10_w8, c1_n10_w9, c1_n10_w10, c1_n10_w11, c1_n10_w12, c1_n10_w13, c1_n10_w14, c1_n10_w15, c1_n10_w16, c1_n10_w17, c1_n10_w18, c1_n10_w19, c1_n10_w20, c1_n10_w21, c1_n10_w22, c1_n10_w23, c1_n10_w24, c1_n10_w25, c1_n10_w26, c1_n10_w27, c1_n10_w28, c1_n10_w29, c1_n10_w30, c1_n10_w31, c1_n10_w32, c1_n10_w33, c1_n10_w34, c1_n10_w35, c1_n10_w36, c1_n10_w37, c1_n10_w38, c1_n10_w39, c1_n10_w40, c1_n10_w41, c1_n10_w42, c1_n10_w43, c1_n10_w44, c1_n10_w45, c1_n10_w46, c1_n10_w47, c1_n10_w48, c1_n10_w49, c1_n10_w50, c1_n10_w51, c1_n10_w52, c1_n10_w53, c1_n10_w54, c1_n10_w55, c1_n10_w56, c1_n10_w57, c1_n10_w58, c1_n10_w59, c1_n10_w60, c1_n10_w61, c1_n10_w62, c1_n10_w63, c1_n10_w64, c1_n10_w65, c1_n10_w66, c1_n10_w67, c1_n10_w68, c1_n10_w69, c1_n10_w70, c1_n10_w71, c1_n10_w72, c1_n10_w73, c1_n10_w74, c1_n10_w75, c1_n10_w76, c1_n10_w77, c1_n10_w78, c1_n10_w79, c1_n10_w80, c1_n10_w81, c1_n10_w82, c1_n10_w83, c1_n10_w84, c1_n10_w85, c1_n10_w86, c1_n10_w87, c1_n10_w88, c1_n10_w89, c1_n10_w90, c1_n10_w91, c1_n10_w92, c1_n10_w93, c1_n10_w94, c1_n10_w95, c1_n10_w96, c1_n10_w97, c1_n10_w98, c1_n10_w99, c1_n10_w100, c1_n11_w1, c1_n11_w2, c1_n11_w3, c1_n11_w4, c1_n11_w5, c1_n11_w6, c1_n11_w7, c1_n11_w8, c1_n11_w9, c1_n11_w10, c1_n11_w11, c1_n11_w12, c1_n11_w13, c1_n11_w14, c1_n11_w15, c1_n11_w16, c1_n11_w17, c1_n11_w18, c1_n11_w19, c1_n11_w20, c1_n11_w21, c1_n11_w22, c1_n11_w23, c1_n11_w24, c1_n11_w25, c1_n11_w26, c1_n11_w27, c1_n11_w28, c1_n11_w29, c1_n11_w30, c1_n11_w31, c1_n11_w32, c1_n11_w33, c1_n11_w34, c1_n11_w35, c1_n11_w36, c1_n11_w37, c1_n11_w38, c1_n11_w39, c1_n11_w40, c1_n11_w41, c1_n11_w42, c1_n11_w43, c1_n11_w44, c1_n11_w45, c1_n11_w46, c1_n11_w47, c1_n11_w48, c1_n11_w49, c1_n11_w50, c1_n11_w51, c1_n11_w52, c1_n11_w53, c1_n11_w54, c1_n11_w55, c1_n11_w56, c1_n11_w57, c1_n11_w58, c1_n11_w59, c1_n11_w60, c1_n11_w61, c1_n11_w62, c1_n11_w63, c1_n11_w64, c1_n11_w65, c1_n11_w66, c1_n11_w67, c1_n11_w68, c1_n11_w69, c1_n11_w70, c1_n11_w71, c1_n11_w72, c1_n11_w73, c1_n11_w74, c1_n11_w75, c1_n11_w76, c1_n11_w77, c1_n11_w78, c1_n11_w79, c1_n11_w80, c1_n11_w81, c1_n11_w82, c1_n11_w83, c1_n11_w84, c1_n11_w85, c1_n11_w86, c1_n11_w87, c1_n11_w88, c1_n11_w89, c1_n11_w90, c1_n11_w91, c1_n11_w92, c1_n11_w93, c1_n11_w94, c1_n11_w95, c1_n11_w96, c1_n11_w97, c1_n11_w98, c1_n11_w99, c1_n11_w100, c1_n12_w1, c1_n12_w2, c1_n12_w3, c1_n12_w4, c1_n12_w5, c1_n12_w6, c1_n12_w7, c1_n12_w8, c1_n12_w9, c1_n12_w10, c1_n12_w11, c1_n12_w12, c1_n12_w13, c1_n12_w14, c1_n12_w15, c1_n12_w16, c1_n12_w17, c1_n12_w18, c1_n12_w19, c1_n12_w20, c1_n12_w21, c1_n12_w22, c1_n12_w23, c1_n12_w24, c1_n12_w25, c1_n12_w26, c1_n12_w27, c1_n12_w28, c1_n12_w29, c1_n12_w30, c1_n12_w31, c1_n12_w32, c1_n12_w33, c1_n12_w34, c1_n12_w35, c1_n12_w36, c1_n12_w37, c1_n12_w38, c1_n12_w39, c1_n12_w40, c1_n12_w41, c1_n12_w42, c1_n12_w43, c1_n12_w44, c1_n12_w45, c1_n12_w46, c1_n12_w47, c1_n12_w48, c1_n12_w49, c1_n12_w50, c1_n12_w51, c1_n12_w52, c1_n12_w53, c1_n12_w54, c1_n12_w55, c1_n12_w56, c1_n12_w57, c1_n12_w58, c1_n12_w59, c1_n12_w60, c1_n12_w61, c1_n12_w62, c1_n12_w63, c1_n12_w64, c1_n12_w65, c1_n12_w66, c1_n12_w67, c1_n12_w68, c1_n12_w69, c1_n12_w70, c1_n12_w71, c1_n12_w72, c1_n12_w73, c1_n12_w74, c1_n12_w75, c1_n12_w76, c1_n12_w77, c1_n12_w78, c1_n12_w79, c1_n12_w80, c1_n12_w81, c1_n12_w82, c1_n12_w83, c1_n12_w84, c1_n12_w85, c1_n12_w86, c1_n12_w87, c1_n12_w88, c1_n12_w89, c1_n12_w90, c1_n12_w91, c1_n12_w92, c1_n12_w93, c1_n12_w94, c1_n12_w95, c1_n12_w96, c1_n12_w97, c1_n12_w98, c1_n12_w99, c1_n12_w100, c1_n13_w1, c1_n13_w2, c1_n13_w3, c1_n13_w4, c1_n13_w5, c1_n13_w6, c1_n13_w7, c1_n13_w8, c1_n13_w9, c1_n13_w10, c1_n13_w11, c1_n13_w12, c1_n13_w13, c1_n13_w14, c1_n13_w15, c1_n13_w16, c1_n13_w17, c1_n13_w18, c1_n13_w19, c1_n13_w20, c1_n13_w21, c1_n13_w22, c1_n13_w23, c1_n13_w24, c1_n13_w25, c1_n13_w26, c1_n13_w27, c1_n13_w28, c1_n13_w29, c1_n13_w30, c1_n13_w31, c1_n13_w32, c1_n13_w33, c1_n13_w34, c1_n13_w35, c1_n13_w36, c1_n13_w37, c1_n13_w38, c1_n13_w39, c1_n13_w40, c1_n13_w41, c1_n13_w42, c1_n13_w43, c1_n13_w44, c1_n13_w45, c1_n13_w46, c1_n13_w47, c1_n13_w48, c1_n13_w49, c1_n13_w50, c1_n13_w51, c1_n13_w52, c1_n13_w53, c1_n13_w54, c1_n13_w55, c1_n13_w56, c1_n13_w57, c1_n13_w58, c1_n13_w59, c1_n13_w60, c1_n13_w61, c1_n13_w62, c1_n13_w63, c1_n13_w64, c1_n13_w65, c1_n13_w66, c1_n13_w67, c1_n13_w68, c1_n13_w69, c1_n13_w70, c1_n13_w71, c1_n13_w72, c1_n13_w73, c1_n13_w74, c1_n13_w75, c1_n13_w76, c1_n13_w77, c1_n13_w78, c1_n13_w79, c1_n13_w80, c1_n13_w81, c1_n13_w82, c1_n13_w83, c1_n13_w84, c1_n13_w85, c1_n13_w86, c1_n13_w87, c1_n13_w88, c1_n13_w89, c1_n13_w90, c1_n13_w91, c1_n13_w92, c1_n13_w93, c1_n13_w94, c1_n13_w95, c1_n13_w96, c1_n13_w97, c1_n13_w98, c1_n13_w99, c1_n13_w100, c1_n14_w1, c1_n14_w2, c1_n14_w3, c1_n14_w4, c1_n14_w5, c1_n14_w6, c1_n14_w7, c1_n14_w8, c1_n14_w9, c1_n14_w10, c1_n14_w11, c1_n14_w12, c1_n14_w13, c1_n14_w14, c1_n14_w15, c1_n14_w16, c1_n14_w17, c1_n14_w18, c1_n14_w19, c1_n14_w20, c1_n14_w21, c1_n14_w22, c1_n14_w23, c1_n14_w24, c1_n14_w25, c1_n14_w26, c1_n14_w27, c1_n14_w28, c1_n14_w29, c1_n14_w30, c1_n14_w31, c1_n14_w32, c1_n14_w33, c1_n14_w34, c1_n14_w35, c1_n14_w36, c1_n14_w37, c1_n14_w38, c1_n14_w39, c1_n14_w40, c1_n14_w41, c1_n14_w42, c1_n14_w43, c1_n14_w44, c1_n14_w45, c1_n14_w46, c1_n14_w47, c1_n14_w48, c1_n14_w49, c1_n14_w50, c1_n14_w51, c1_n14_w52, c1_n14_w53, c1_n14_w54, c1_n14_w55, c1_n14_w56, c1_n14_w57, c1_n14_w58, c1_n14_w59, c1_n14_w60, c1_n14_w61, c1_n14_w62, c1_n14_w63, c1_n14_w64, c1_n14_w65, c1_n14_w66, c1_n14_w67, c1_n14_w68, c1_n14_w69, c1_n14_w70, c1_n14_w71, c1_n14_w72, c1_n14_w73, c1_n14_w74, c1_n14_w75, c1_n14_w76, c1_n14_w77, c1_n14_w78, c1_n14_w79, c1_n14_w80, c1_n14_w81, c1_n14_w82, c1_n14_w83, c1_n14_w84, c1_n14_w85, c1_n14_w86, c1_n14_w87, c1_n14_w88, c1_n14_w89, c1_n14_w90, c1_n14_w91, c1_n14_w92, c1_n14_w93, c1_n14_w94, c1_n14_w95, c1_n14_w96, c1_n14_w97, c1_n14_w98, c1_n14_w99, c1_n14_w100, c1_n15_w1, c1_n15_w2, c1_n15_w3, c1_n15_w4, c1_n15_w5, c1_n15_w6, c1_n15_w7, c1_n15_w8, c1_n15_w9, c1_n15_w10, c1_n15_w11, c1_n15_w12, c1_n15_w13, c1_n15_w14, c1_n15_w15, c1_n15_w16, c1_n15_w17, c1_n15_w18, c1_n15_w19, c1_n15_w20, c1_n15_w21, c1_n15_w22, c1_n15_w23, c1_n15_w24, c1_n15_w25, c1_n15_w26, c1_n15_w27, c1_n15_w28, c1_n15_w29, c1_n15_w30, c1_n15_w31, c1_n15_w32, c1_n15_w33, c1_n15_w34, c1_n15_w35, c1_n15_w36, c1_n15_w37, c1_n15_w38, c1_n15_w39, c1_n15_w40, c1_n15_w41, c1_n15_w42, c1_n15_w43, c1_n15_w44, c1_n15_w45, c1_n15_w46, c1_n15_w47, c1_n15_w48, c1_n15_w49, c1_n15_w50, c1_n15_w51, c1_n15_w52, c1_n15_w53, c1_n15_w54, c1_n15_w55, c1_n15_w56, c1_n15_w57, c1_n15_w58, c1_n15_w59, c1_n15_w60, c1_n15_w61, c1_n15_w62, c1_n15_w63, c1_n15_w64, c1_n15_w65, c1_n15_w66, c1_n15_w67, c1_n15_w68, c1_n15_w69, c1_n15_w70, c1_n15_w71, c1_n15_w72, c1_n15_w73, c1_n15_w74, c1_n15_w75, c1_n15_w76, c1_n15_w77, c1_n15_w78, c1_n15_w79, c1_n15_w80, c1_n15_w81, c1_n15_w82, c1_n15_w83, c1_n15_w84, c1_n15_w85, c1_n15_w86, c1_n15_w87, c1_n15_w88, c1_n15_w89, c1_n15_w90, c1_n15_w91, c1_n15_w92, c1_n15_w93, c1_n15_w94, c1_n15_w95, c1_n15_w96, c1_n15_w97, c1_n15_w98, c1_n15_w99, c1_n15_w100, c1_n16_w1, c1_n16_w2, c1_n16_w3, c1_n16_w4, c1_n16_w5, c1_n16_w6, c1_n16_w7, c1_n16_w8, c1_n16_w9, c1_n16_w10, c1_n16_w11, c1_n16_w12, c1_n16_w13, c1_n16_w14, c1_n16_w15, c1_n16_w16, c1_n16_w17, c1_n16_w18, c1_n16_w19, c1_n16_w20, c1_n16_w21, c1_n16_w22, c1_n16_w23, c1_n16_w24, c1_n16_w25, c1_n16_w26, c1_n16_w27, c1_n16_w28, c1_n16_w29, c1_n16_w30, c1_n16_w31, c1_n16_w32, c1_n16_w33, c1_n16_w34, c1_n16_w35, c1_n16_w36, c1_n16_w37, c1_n16_w38, c1_n16_w39, c1_n16_w40, c1_n16_w41, c1_n16_w42, c1_n16_w43, c1_n16_w44, c1_n16_w45, c1_n16_w46, c1_n16_w47, c1_n16_w48, c1_n16_w49, c1_n16_w50, c1_n16_w51, c1_n16_w52, c1_n16_w53, c1_n16_w54, c1_n16_w55, c1_n16_w56, c1_n16_w57, c1_n16_w58, c1_n16_w59, c1_n16_w60, c1_n16_w61, c1_n16_w62, c1_n16_w63, c1_n16_w64, c1_n16_w65, c1_n16_w66, c1_n16_w67, c1_n16_w68, c1_n16_w69, c1_n16_w70, c1_n16_w71, c1_n16_w72, c1_n16_w73, c1_n16_w74, c1_n16_w75, c1_n16_w76, c1_n16_w77, c1_n16_w78, c1_n16_w79, c1_n16_w80, c1_n16_w81, c1_n16_w82, c1_n16_w83, c1_n16_w84, c1_n16_w85, c1_n16_w86, c1_n16_w87, c1_n16_w88, c1_n16_w89, c1_n16_w90, c1_n16_w91, c1_n16_w92, c1_n16_w93, c1_n16_w94, c1_n16_w95, c1_n16_w96, c1_n16_w97, c1_n16_w98, c1_n16_w99, c1_n16_w100, c1_n17_w1, c1_n17_w2, c1_n17_w3, c1_n17_w4, c1_n17_w5, c1_n17_w6, c1_n17_w7, c1_n17_w8, c1_n17_w9, c1_n17_w10, c1_n17_w11, c1_n17_w12, c1_n17_w13, c1_n17_w14, c1_n17_w15, c1_n17_w16, c1_n17_w17, c1_n17_w18, c1_n17_w19, c1_n17_w20, c1_n17_w21, c1_n17_w22, c1_n17_w23, c1_n17_w24, c1_n17_w25, c1_n17_w26, c1_n17_w27, c1_n17_w28, c1_n17_w29, c1_n17_w30, c1_n17_w31, c1_n17_w32, c1_n17_w33, c1_n17_w34, c1_n17_w35, c1_n17_w36, c1_n17_w37, c1_n17_w38, c1_n17_w39, c1_n17_w40, c1_n17_w41, c1_n17_w42, c1_n17_w43, c1_n17_w44, c1_n17_w45, c1_n17_w46, c1_n17_w47, c1_n17_w48, c1_n17_w49, c1_n17_w50, c1_n17_w51, c1_n17_w52, c1_n17_w53, c1_n17_w54, c1_n17_w55, c1_n17_w56, c1_n17_w57, c1_n17_w58, c1_n17_w59, c1_n17_w60, c1_n17_w61, c1_n17_w62, c1_n17_w63, c1_n17_w64, c1_n17_w65, c1_n17_w66, c1_n17_w67, c1_n17_w68, c1_n17_w69, c1_n17_w70, c1_n17_w71, c1_n17_w72, c1_n17_w73, c1_n17_w74, c1_n17_w75, c1_n17_w76, c1_n17_w77, c1_n17_w78, c1_n17_w79, c1_n17_w80, c1_n17_w81, c1_n17_w82, c1_n17_w83, c1_n17_w84, c1_n17_w85, c1_n17_w86, c1_n17_w87, c1_n17_w88, c1_n17_w89, c1_n17_w90, c1_n17_w91, c1_n17_w92, c1_n17_w93, c1_n17_w94, c1_n17_w95, c1_n17_w96, c1_n17_w97, c1_n17_w98, c1_n17_w99, c1_n17_w100, c1_n18_w1, c1_n18_w2, c1_n18_w3, c1_n18_w4, c1_n18_w5, c1_n18_w6, c1_n18_w7, c1_n18_w8, c1_n18_w9, c1_n18_w10, c1_n18_w11, c1_n18_w12, c1_n18_w13, c1_n18_w14, c1_n18_w15, c1_n18_w16, c1_n18_w17, c1_n18_w18, c1_n18_w19, c1_n18_w20, c1_n18_w21, c1_n18_w22, c1_n18_w23, c1_n18_w24, c1_n18_w25, c1_n18_w26, c1_n18_w27, c1_n18_w28, c1_n18_w29, c1_n18_w30, c1_n18_w31, c1_n18_w32, c1_n18_w33, c1_n18_w34, c1_n18_w35, c1_n18_w36, c1_n18_w37, c1_n18_w38, c1_n18_w39, c1_n18_w40, c1_n18_w41, c1_n18_w42, c1_n18_w43, c1_n18_w44, c1_n18_w45, c1_n18_w46, c1_n18_w47, c1_n18_w48, c1_n18_w49, c1_n18_w50, c1_n18_w51, c1_n18_w52, c1_n18_w53, c1_n18_w54, c1_n18_w55, c1_n18_w56, c1_n18_w57, c1_n18_w58, c1_n18_w59, c1_n18_w60, c1_n18_w61, c1_n18_w62, c1_n18_w63, c1_n18_w64, c1_n18_w65, c1_n18_w66, c1_n18_w67, c1_n18_w68, c1_n18_w69, c1_n18_w70, c1_n18_w71, c1_n18_w72, c1_n18_w73, c1_n18_w74, c1_n18_w75, c1_n18_w76, c1_n18_w77, c1_n18_w78, c1_n18_w79, c1_n18_w80, c1_n18_w81, c1_n18_w82, c1_n18_w83, c1_n18_w84, c1_n18_w85, c1_n18_w86, c1_n18_w87, c1_n18_w88, c1_n18_w89, c1_n18_w90, c1_n18_w91, c1_n18_w92, c1_n18_w93, c1_n18_w94, c1_n18_w95, c1_n18_w96, c1_n18_w97, c1_n18_w98, c1_n18_w99, c1_n18_w100, c1_n19_w1, c1_n19_w2, c1_n19_w3, c1_n19_w4, c1_n19_w5, c1_n19_w6, c1_n19_w7, c1_n19_w8, c1_n19_w9, c1_n19_w10, c1_n19_w11, c1_n19_w12, c1_n19_w13, c1_n19_w14, c1_n19_w15, c1_n19_w16, c1_n19_w17, c1_n19_w18, c1_n19_w19, c1_n19_w20, c1_n19_w21, c1_n19_w22, c1_n19_w23, c1_n19_w24, c1_n19_w25, c1_n19_w26, c1_n19_w27, c1_n19_w28, c1_n19_w29, c1_n19_w30, c1_n19_w31, c1_n19_w32, c1_n19_w33, c1_n19_w34, c1_n19_w35, c1_n19_w36, c1_n19_w37, c1_n19_w38, c1_n19_w39, c1_n19_w40, c1_n19_w41, c1_n19_w42, c1_n19_w43, c1_n19_w44, c1_n19_w45, c1_n19_w46, c1_n19_w47, c1_n19_w48, c1_n19_w49, c1_n19_w50, c1_n19_w51, c1_n19_w52, c1_n19_w53, c1_n19_w54, c1_n19_w55, c1_n19_w56, c1_n19_w57, c1_n19_w58, c1_n19_w59, c1_n19_w60, c1_n19_w61, c1_n19_w62, c1_n19_w63, c1_n19_w64, c1_n19_w65, c1_n19_w66, c1_n19_w67, c1_n19_w68, c1_n19_w69, c1_n19_w70, c1_n19_w71, c1_n19_w72, c1_n19_w73, c1_n19_w74, c1_n19_w75, c1_n19_w76, c1_n19_w77, c1_n19_w78, c1_n19_w79, c1_n19_w80, c1_n19_w81, c1_n19_w82, c1_n19_w83, c1_n19_w84, c1_n19_w85, c1_n19_w86, c1_n19_w87, c1_n19_w88, c1_n19_w89, c1_n19_w90, c1_n19_w91, c1_n19_w92, c1_n19_w93, c1_n19_w94, c1_n19_w95, c1_n19_w96, c1_n19_w97, c1_n19_w98, c1_n19_w99, c1_n19_w100, c1_n20_w1, c1_n20_w2, c1_n20_w3, c1_n20_w4, c1_n20_w5, c1_n20_w6, c1_n20_w7, c1_n20_w8, c1_n20_w9, c1_n20_w10, c1_n20_w11, c1_n20_w12, c1_n20_w13, c1_n20_w14, c1_n20_w15, c1_n20_w16, c1_n20_w17, c1_n20_w18, c1_n20_w19, c1_n20_w20, c1_n20_w21, c1_n20_w22, c1_n20_w23, c1_n20_w24, c1_n20_w25, c1_n20_w26, c1_n20_w27, c1_n20_w28, c1_n20_w29, c1_n20_w30, c1_n20_w31, c1_n20_w32, c1_n20_w33, c1_n20_w34, c1_n20_w35, c1_n20_w36, c1_n20_w37, c1_n20_w38, c1_n20_w39, c1_n20_w40, c1_n20_w41, c1_n20_w42, c1_n20_w43, c1_n20_w44, c1_n20_w45, c1_n20_w46, c1_n20_w47, c1_n20_w48, c1_n20_w49, c1_n20_w50, c1_n20_w51, c1_n20_w52, c1_n20_w53, c1_n20_w54, c1_n20_w55, c1_n20_w56, c1_n20_w57, c1_n20_w58, c1_n20_w59, c1_n20_w60, c1_n20_w61, c1_n20_w62, c1_n20_w63, c1_n20_w64, c1_n20_w65, c1_n20_w66, c1_n20_w67, c1_n20_w68, c1_n20_w69, c1_n20_w70, c1_n20_w71, c1_n20_w72, c1_n20_w73, c1_n20_w74, c1_n20_w75, c1_n20_w76, c1_n20_w77, c1_n20_w78, c1_n20_w79, c1_n20_w80, c1_n20_w81, c1_n20_w82, c1_n20_w83, c1_n20_w84, c1_n20_w85, c1_n20_w86, c1_n20_w87, c1_n20_w88, c1_n20_w89, c1_n20_w90, c1_n20_w91, c1_n20_w92, c1_n20_w93, c1_n20_w94, c1_n20_w95, c1_n20_w96, c1_n20_w97, c1_n20_w98, c1_n20_w99, c1_n20_w100, c1_n21_w1, c1_n21_w2, c1_n21_w3, c1_n21_w4, c1_n21_w5, c1_n21_w6, c1_n21_w7, c1_n21_w8, c1_n21_w9, c1_n21_w10, c1_n21_w11, c1_n21_w12, c1_n21_w13, c1_n21_w14, c1_n21_w15, c1_n21_w16, c1_n21_w17, c1_n21_w18, c1_n21_w19, c1_n21_w20, c1_n21_w21, c1_n21_w22, c1_n21_w23, c1_n21_w24, c1_n21_w25, c1_n21_w26, c1_n21_w27, c1_n21_w28, c1_n21_w29, c1_n21_w30, c1_n21_w31, c1_n21_w32, c1_n21_w33, c1_n21_w34, c1_n21_w35, c1_n21_w36, c1_n21_w37, c1_n21_w38, c1_n21_w39, c1_n21_w40, c1_n21_w41, c1_n21_w42, c1_n21_w43, c1_n21_w44, c1_n21_w45, c1_n21_w46, c1_n21_w47, c1_n21_w48, c1_n21_w49, c1_n21_w50, c1_n21_w51, c1_n21_w52, c1_n21_w53, c1_n21_w54, c1_n21_w55, c1_n21_w56, c1_n21_w57, c1_n21_w58, c1_n21_w59, c1_n21_w60, c1_n21_w61, c1_n21_w62, c1_n21_w63, c1_n21_w64, c1_n21_w65, c1_n21_w66, c1_n21_w67, c1_n21_w68, c1_n21_w69, c1_n21_w70, c1_n21_w71, c1_n21_w72, c1_n21_w73, c1_n21_w74, c1_n21_w75, c1_n21_w76, c1_n21_w77, c1_n21_w78, c1_n21_w79, c1_n21_w80, c1_n21_w81, c1_n21_w82, c1_n21_w83, c1_n21_w84, c1_n21_w85, c1_n21_w86, c1_n21_w87, c1_n21_w88, c1_n21_w89, c1_n21_w90, c1_n21_w91, c1_n21_w92, c1_n21_w93, c1_n21_w94, c1_n21_w95, c1_n21_w96, c1_n21_w97, c1_n21_w98, c1_n21_w99, c1_n21_w100, c1_n22_w1, c1_n22_w2, c1_n22_w3, c1_n22_w4, c1_n22_w5, c1_n22_w6, c1_n22_w7, c1_n22_w8, c1_n22_w9, c1_n22_w10, c1_n22_w11, c1_n22_w12, c1_n22_w13, c1_n22_w14, c1_n22_w15, c1_n22_w16, c1_n22_w17, c1_n22_w18, c1_n22_w19, c1_n22_w20, c1_n22_w21, c1_n22_w22, c1_n22_w23, c1_n22_w24, c1_n22_w25, c1_n22_w26, c1_n22_w27, c1_n22_w28, c1_n22_w29, c1_n22_w30, c1_n22_w31, c1_n22_w32, c1_n22_w33, c1_n22_w34, c1_n22_w35, c1_n22_w36, c1_n22_w37, c1_n22_w38, c1_n22_w39, c1_n22_w40, c1_n22_w41, c1_n22_w42, c1_n22_w43, c1_n22_w44, c1_n22_w45, c1_n22_w46, c1_n22_w47, c1_n22_w48, c1_n22_w49, c1_n22_w50, c1_n22_w51, c1_n22_w52, c1_n22_w53, c1_n22_w54, c1_n22_w55, c1_n22_w56, c1_n22_w57, c1_n22_w58, c1_n22_w59, c1_n22_w60, c1_n22_w61, c1_n22_w62, c1_n22_w63, c1_n22_w64, c1_n22_w65, c1_n22_w66, c1_n22_w67, c1_n22_w68, c1_n22_w69, c1_n22_w70, c1_n22_w71, c1_n22_w72, c1_n22_w73, c1_n22_w74, c1_n22_w75, c1_n22_w76, c1_n22_w77, c1_n22_w78, c1_n22_w79, c1_n22_w80, c1_n22_w81, c1_n22_w82, c1_n22_w83, c1_n22_w84, c1_n22_w85, c1_n22_w86, c1_n22_w87, c1_n22_w88, c1_n22_w89, c1_n22_w90, c1_n22_w91, c1_n22_w92, c1_n22_w93, c1_n22_w94, c1_n22_w95, c1_n22_w96, c1_n22_w97, c1_n22_w98, c1_n22_w99, c1_n22_w100, c1_n23_w1, c1_n23_w2, c1_n23_w3, c1_n23_w4, c1_n23_w5, c1_n23_w6, c1_n23_w7, c1_n23_w8, c1_n23_w9, c1_n23_w10, c1_n23_w11, c1_n23_w12, c1_n23_w13, c1_n23_w14, c1_n23_w15, c1_n23_w16, c1_n23_w17, c1_n23_w18, c1_n23_w19, c1_n23_w20, c1_n23_w21, c1_n23_w22, c1_n23_w23, c1_n23_w24, c1_n23_w25, c1_n23_w26, c1_n23_w27, c1_n23_w28, c1_n23_w29, c1_n23_w30, c1_n23_w31, c1_n23_w32, c1_n23_w33, c1_n23_w34, c1_n23_w35, c1_n23_w36, c1_n23_w37, c1_n23_w38, c1_n23_w39, c1_n23_w40, c1_n23_w41, c1_n23_w42, c1_n23_w43, c1_n23_w44, c1_n23_w45, c1_n23_w46, c1_n23_w47, c1_n23_w48, c1_n23_w49, c1_n23_w50, c1_n23_w51, c1_n23_w52, c1_n23_w53, c1_n23_w54, c1_n23_w55, c1_n23_w56, c1_n23_w57, c1_n23_w58, c1_n23_w59, c1_n23_w60, c1_n23_w61, c1_n23_w62, c1_n23_w63, c1_n23_w64, c1_n23_w65, c1_n23_w66, c1_n23_w67, c1_n23_w68, c1_n23_w69, c1_n23_w70, c1_n23_w71, c1_n23_w72, c1_n23_w73, c1_n23_w74, c1_n23_w75, c1_n23_w76, c1_n23_w77, c1_n23_w78, c1_n23_w79, c1_n23_w80, c1_n23_w81, c1_n23_w82, c1_n23_w83, c1_n23_w84, c1_n23_w85, c1_n23_w86, c1_n23_w87, c1_n23_w88, c1_n23_w89, c1_n23_w90, c1_n23_w91, c1_n23_w92, c1_n23_w93, c1_n23_w94, c1_n23_w95, c1_n23_w96, c1_n23_w97, c1_n23_w98, c1_n23_w99, c1_n23_w100, c1_n24_w1, c1_n24_w2, c1_n24_w3, c1_n24_w4, c1_n24_w5, c1_n24_w6, c1_n24_w7, c1_n24_w8, c1_n24_w9, c1_n24_w10, c1_n24_w11, c1_n24_w12, c1_n24_w13, c1_n24_w14, c1_n24_w15, c1_n24_w16, c1_n24_w17, c1_n24_w18, c1_n24_w19, c1_n24_w20, c1_n24_w21, c1_n24_w22, c1_n24_w23, c1_n24_w24, c1_n24_w25, c1_n24_w26, c1_n24_w27, c1_n24_w28, c1_n24_w29, c1_n24_w30, c1_n24_w31, c1_n24_w32, c1_n24_w33, c1_n24_w34, c1_n24_w35, c1_n24_w36, c1_n24_w37, c1_n24_w38, c1_n24_w39, c1_n24_w40, c1_n24_w41, c1_n24_w42, c1_n24_w43, c1_n24_w44, c1_n24_w45, c1_n24_w46, c1_n24_w47, c1_n24_w48, c1_n24_w49, c1_n24_w50, c1_n24_w51, c1_n24_w52, c1_n24_w53, c1_n24_w54, c1_n24_w55, c1_n24_w56, c1_n24_w57, c1_n24_w58, c1_n24_w59, c1_n24_w60, c1_n24_w61, c1_n24_w62, c1_n24_w63, c1_n24_w64, c1_n24_w65, c1_n24_w66, c1_n24_w67, c1_n24_w68, c1_n24_w69, c1_n24_w70, c1_n24_w71, c1_n24_w72, c1_n24_w73, c1_n24_w74, c1_n24_w75, c1_n24_w76, c1_n24_w77, c1_n24_w78, c1_n24_w79, c1_n24_w80, c1_n24_w81, c1_n24_w82, c1_n24_w83, c1_n24_w84, c1_n24_w85, c1_n24_w86, c1_n24_w87, c1_n24_w88, c1_n24_w89, c1_n24_w90, c1_n24_w91, c1_n24_w92, c1_n24_w93, c1_n24_w94, c1_n24_w95, c1_n24_w96, c1_n24_w97, c1_n24_w98, c1_n24_w99, c1_n24_w100, c1_n25_w1, c1_n25_w2, c1_n25_w3, c1_n25_w4, c1_n25_w5, c1_n25_w6, c1_n25_w7, c1_n25_w8, c1_n25_w9, c1_n25_w10, c1_n25_w11, c1_n25_w12, c1_n25_w13, c1_n25_w14, c1_n25_w15, c1_n25_w16, c1_n25_w17, c1_n25_w18, c1_n25_w19, c1_n25_w20, c1_n25_w21, c1_n25_w22, c1_n25_w23, c1_n25_w24, c1_n25_w25, c1_n25_w26, c1_n25_w27, c1_n25_w28, c1_n25_w29, c1_n25_w30, c1_n25_w31, c1_n25_w32, c1_n25_w33, c1_n25_w34, c1_n25_w35, c1_n25_w36, c1_n25_w37, c1_n25_w38, c1_n25_w39, c1_n25_w40, c1_n25_w41, c1_n25_w42, c1_n25_w43, c1_n25_w44, c1_n25_w45, c1_n25_w46, c1_n25_w47, c1_n25_w48, c1_n25_w49, c1_n25_w50, c1_n25_w51, c1_n25_w52, c1_n25_w53, c1_n25_w54, c1_n25_w55, c1_n25_w56, c1_n25_w57, c1_n25_w58, c1_n25_w59, c1_n25_w60, c1_n25_w61, c1_n25_w62, c1_n25_w63, c1_n25_w64, c1_n25_w65, c1_n25_w66, c1_n25_w67, c1_n25_w68, c1_n25_w69, c1_n25_w70, c1_n25_w71, c1_n25_w72, c1_n25_w73, c1_n25_w74, c1_n25_w75, c1_n25_w76, c1_n25_w77, c1_n25_w78, c1_n25_w79, c1_n25_w80, c1_n25_w81, c1_n25_w82, c1_n25_w83, c1_n25_w84, c1_n25_w85, c1_n25_w86, c1_n25_w87, c1_n25_w88, c1_n25_w89, c1_n25_w90, c1_n25_w91, c1_n25_w92, c1_n25_w93, c1_n25_w94, c1_n25_w95, c1_n25_w96, c1_n25_w97, c1_n25_w98, c1_n25_w99, c1_n25_w100, c1_n26_w1, c1_n26_w2, c1_n26_w3, c1_n26_w4, c1_n26_w5, c1_n26_w6, c1_n26_w7, c1_n26_w8, c1_n26_w9, c1_n26_w10, c1_n26_w11, c1_n26_w12, c1_n26_w13, c1_n26_w14, c1_n26_w15, c1_n26_w16, c1_n26_w17, c1_n26_w18, c1_n26_w19, c1_n26_w20, c1_n26_w21, c1_n26_w22, c1_n26_w23, c1_n26_w24, c1_n26_w25, c1_n26_w26, c1_n26_w27, c1_n26_w28, c1_n26_w29, c1_n26_w30, c1_n26_w31, c1_n26_w32, c1_n26_w33, c1_n26_w34, c1_n26_w35, c1_n26_w36, c1_n26_w37, c1_n26_w38, c1_n26_w39, c1_n26_w40, c1_n26_w41, c1_n26_w42, c1_n26_w43, c1_n26_w44, c1_n26_w45, c1_n26_w46, c1_n26_w47, c1_n26_w48, c1_n26_w49, c1_n26_w50, c1_n26_w51, c1_n26_w52, c1_n26_w53, c1_n26_w54, c1_n26_w55, c1_n26_w56, c1_n26_w57, c1_n26_w58, c1_n26_w59, c1_n26_w60, c1_n26_w61, c1_n26_w62, c1_n26_w63, c1_n26_w64, c1_n26_w65, c1_n26_w66, c1_n26_w67, c1_n26_w68, c1_n26_w69, c1_n26_w70, c1_n26_w71, c1_n26_w72, c1_n26_w73, c1_n26_w74, c1_n26_w75, c1_n26_w76, c1_n26_w77, c1_n26_w78, c1_n26_w79, c1_n26_w80, c1_n26_w81, c1_n26_w82, c1_n26_w83, c1_n26_w84, c1_n26_w85, c1_n26_w86, c1_n26_w87, c1_n26_w88, c1_n26_w89, c1_n26_w90, c1_n26_w91, c1_n26_w92, c1_n26_w93, c1_n26_w94, c1_n26_w95, c1_n26_w96, c1_n26_w97, c1_n26_w98, c1_n26_w99, c1_n26_w100, c1_n27_w1, c1_n27_w2, c1_n27_w3, c1_n27_w4, c1_n27_w5, c1_n27_w6, c1_n27_w7, c1_n27_w8, c1_n27_w9, c1_n27_w10, c1_n27_w11, c1_n27_w12, c1_n27_w13, c1_n27_w14, c1_n27_w15, c1_n27_w16, c1_n27_w17, c1_n27_w18, c1_n27_w19, c1_n27_w20, c1_n27_w21, c1_n27_w22, c1_n27_w23, c1_n27_w24, c1_n27_w25, c1_n27_w26, c1_n27_w27, c1_n27_w28, c1_n27_w29, c1_n27_w30, c1_n27_w31, c1_n27_w32, c1_n27_w33, c1_n27_w34, c1_n27_w35, c1_n27_w36, c1_n27_w37, c1_n27_w38, c1_n27_w39, c1_n27_w40, c1_n27_w41, c1_n27_w42, c1_n27_w43, c1_n27_w44, c1_n27_w45, c1_n27_w46, c1_n27_w47, c1_n27_w48, c1_n27_w49, c1_n27_w50, c1_n27_w51, c1_n27_w52, c1_n27_w53, c1_n27_w54, c1_n27_w55, c1_n27_w56, c1_n27_w57, c1_n27_w58, c1_n27_w59, c1_n27_w60, c1_n27_w61, c1_n27_w62, c1_n27_w63, c1_n27_w64, c1_n27_w65, c1_n27_w66, c1_n27_w67, c1_n27_w68, c1_n27_w69, c1_n27_w70, c1_n27_w71, c1_n27_w72, c1_n27_w73, c1_n27_w74, c1_n27_w75, c1_n27_w76, c1_n27_w77, c1_n27_w78, c1_n27_w79, c1_n27_w80, c1_n27_w81, c1_n27_w82, c1_n27_w83, c1_n27_w84, c1_n27_w85, c1_n27_w86, c1_n27_w87, c1_n27_w88, c1_n27_w89, c1_n27_w90, c1_n27_w91, c1_n27_w92, c1_n27_w93, c1_n27_w94, c1_n27_w95, c1_n27_w96, c1_n27_w97, c1_n27_w98, c1_n27_w99, c1_n27_w100, c1_n28_w1, c1_n28_w2, c1_n28_w3, c1_n28_w4, c1_n28_w5, c1_n28_w6, c1_n28_w7, c1_n28_w8, c1_n28_w9, c1_n28_w10, c1_n28_w11, c1_n28_w12, c1_n28_w13, c1_n28_w14, c1_n28_w15, c1_n28_w16, c1_n28_w17, c1_n28_w18, c1_n28_w19, c1_n28_w20, c1_n28_w21, c1_n28_w22, c1_n28_w23, c1_n28_w24, c1_n28_w25, c1_n28_w26, c1_n28_w27, c1_n28_w28, c1_n28_w29, c1_n28_w30, c1_n28_w31, c1_n28_w32, c1_n28_w33, c1_n28_w34, c1_n28_w35, c1_n28_w36, c1_n28_w37, c1_n28_w38, c1_n28_w39, c1_n28_w40, c1_n28_w41, c1_n28_w42, c1_n28_w43, c1_n28_w44, c1_n28_w45, c1_n28_w46, c1_n28_w47, c1_n28_w48, c1_n28_w49, c1_n28_w50, c1_n28_w51, c1_n28_w52, c1_n28_w53, c1_n28_w54, c1_n28_w55, c1_n28_w56, c1_n28_w57, c1_n28_w58, c1_n28_w59, c1_n28_w60, c1_n28_w61, c1_n28_w62, c1_n28_w63, c1_n28_w64, c1_n28_w65, c1_n28_w66, c1_n28_w67, c1_n28_w68, c1_n28_w69, c1_n28_w70, c1_n28_w71, c1_n28_w72, c1_n28_w73, c1_n28_w74, c1_n28_w75, c1_n28_w76, c1_n28_w77, c1_n28_w78, c1_n28_w79, c1_n28_w80, c1_n28_w81, c1_n28_w82, c1_n28_w83, c1_n28_w84, c1_n28_w85, c1_n28_w86, c1_n28_w87, c1_n28_w88, c1_n28_w89, c1_n28_w90, c1_n28_w91, c1_n28_w92, c1_n28_w93, c1_n28_w94, c1_n28_w95, c1_n28_w96, c1_n28_w97, c1_n28_w98, c1_n28_w99, c1_n28_w100, c1_n29_w1, c1_n29_w2, c1_n29_w3, c1_n29_w4, c1_n29_w5, c1_n29_w6, c1_n29_w7, c1_n29_w8, c1_n29_w9, c1_n29_w10, c1_n29_w11, c1_n29_w12, c1_n29_w13, c1_n29_w14, c1_n29_w15, c1_n29_w16, c1_n29_w17, c1_n29_w18, c1_n29_w19, c1_n29_w20, c1_n29_w21, c1_n29_w22, c1_n29_w23, c1_n29_w24, c1_n29_w25, c1_n29_w26, c1_n29_w27, c1_n29_w28, c1_n29_w29, c1_n29_w30, c1_n29_w31, c1_n29_w32, c1_n29_w33, c1_n29_w34, c1_n29_w35, c1_n29_w36, c1_n29_w37, c1_n29_w38, c1_n29_w39, c1_n29_w40, c1_n29_w41, c1_n29_w42, c1_n29_w43, c1_n29_w44, c1_n29_w45, c1_n29_w46, c1_n29_w47, c1_n29_w48, c1_n29_w49, c1_n29_w50, c1_n29_w51, c1_n29_w52, c1_n29_w53, c1_n29_w54, c1_n29_w55, c1_n29_w56, c1_n29_w57, c1_n29_w58, c1_n29_w59, c1_n29_w60, c1_n29_w61, c1_n29_w62, c1_n29_w63, c1_n29_w64, c1_n29_w65, c1_n29_w66, c1_n29_w67, c1_n29_w68, c1_n29_w69, c1_n29_w70, c1_n29_w71, c1_n29_w72, c1_n29_w73, c1_n29_w74, c1_n29_w75, c1_n29_w76, c1_n29_w77, c1_n29_w78, c1_n29_w79, c1_n29_w80, c1_n29_w81, c1_n29_w82, c1_n29_w83, c1_n29_w84, c1_n29_w85, c1_n29_w86, c1_n29_w87, c1_n29_w88, c1_n29_w89, c1_n29_w90, c1_n29_w91, c1_n29_w92, c1_n29_w93, c1_n29_w94, c1_n29_w95, c1_n29_w96, c1_n29_w97, c1_n29_w98, c1_n29_w99, c1_n29_w100: IN signed(7 DOWNTO 0);
    ----------------------------------------------
    c1_n0_y, c1_n1_y, c1_n2_y, c1_n3_y, c1_n4_y, c1_n5_y, c1_n6_y, c1_n7_y, c1_n8_y, c1_n9_y, c1_n10_y, c1_n11_y, c1_n12_y, c1_n13_y, c1_n14_y, c1_n15_y, c1_n16_y, c1_n17_y, c1_n18_y, c1_n19_y, c1_n20_y, c1_n21_y, c1_n22_y, c1_n23_y, c1_n24_y, c1_n25_y, c1_n26_y, c1_n27_y, c1_n28_y, c1_n29_y: OUT signed(7 DOWNTO 0)
    );
end ENTITY;

ARCHITECTURE arch OF  camada1_Leaky_ReLU_30neuron_8bits_100n_signed  IS 
BEGIN

neuron_inst_0: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n0_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n0_w1, 
            w2=> c1_n0_w2, 
            w3=> c1_n0_w3, 
            w4=> c1_n0_w4, 
            w5=> c1_n0_w5, 
            w6=> c1_n0_w6, 
            w7=> c1_n0_w7, 
            w8=> c1_n0_w8, 
            w9=> c1_n0_w9, 
            w10=> c1_n0_w10, 
            w11=> c1_n0_w11, 
            w12=> c1_n0_w12, 
            w13=> c1_n0_w13, 
            w14=> c1_n0_w14, 
            w15=> c1_n0_w15, 
            w16=> c1_n0_w16, 
            w17=> c1_n0_w17, 
            w18=> c1_n0_w18, 
            w19=> c1_n0_w19, 
            w20=> c1_n0_w20, 
            w21=> c1_n0_w21, 
            w22=> c1_n0_w22, 
            w23=> c1_n0_w23, 
            w24=> c1_n0_w24, 
            w25=> c1_n0_w25, 
            w26=> c1_n0_w26, 
            w27=> c1_n0_w27, 
            w28=> c1_n0_w28, 
            w29=> c1_n0_w29, 
            w30=> c1_n0_w30, 
            w31=> c1_n0_w31, 
            w32=> c1_n0_w32, 
            w33=> c1_n0_w33, 
            w34=> c1_n0_w34, 
            w35=> c1_n0_w35, 
            w36=> c1_n0_w36, 
            w37=> c1_n0_w37, 
            w38=> c1_n0_w38, 
            w39=> c1_n0_w39, 
            w40=> c1_n0_w40, 
            w41=> c1_n0_w41, 
            w42=> c1_n0_w42, 
            w43=> c1_n0_w43, 
            w44=> c1_n0_w44, 
            w45=> c1_n0_w45, 
            w46=> c1_n0_w46, 
            w47=> c1_n0_w47, 
            w48=> c1_n0_w48, 
            w49=> c1_n0_w49, 
            w50=> c1_n0_w50, 
            w51=> c1_n0_w51, 
            w52=> c1_n0_w52, 
            w53=> c1_n0_w53, 
            w54=> c1_n0_w54, 
            w55=> c1_n0_w55, 
            w56=> c1_n0_w56, 
            w57=> c1_n0_w57, 
            w58=> c1_n0_w58, 
            w59=> c1_n0_w59, 
            w60=> c1_n0_w60, 
            w61=> c1_n0_w61, 
            w62=> c1_n0_w62, 
            w63=> c1_n0_w63, 
            w64=> c1_n0_w64, 
            w65=> c1_n0_w65, 
            w66=> c1_n0_w66, 
            w67=> c1_n0_w67, 
            w68=> c1_n0_w68, 
            w69=> c1_n0_w69, 
            w70=> c1_n0_w70, 
            w71=> c1_n0_w71, 
            w72=> c1_n0_w72, 
            w73=> c1_n0_w73, 
            w74=> c1_n0_w74, 
            w75=> c1_n0_w75, 
            w76=> c1_n0_w76, 
            w77=> c1_n0_w77, 
            w78=> c1_n0_w78, 
            w79=> c1_n0_w79, 
            w80=> c1_n0_w80, 
            w81=> c1_n0_w81, 
            w82=> c1_n0_w82, 
            w83=> c1_n0_w83, 
            w84=> c1_n0_w84, 
            w85=> c1_n0_w85, 
            w86=> c1_n0_w86, 
            w87=> c1_n0_w87, 
            w88=> c1_n0_w88, 
            w89=> c1_n0_w89, 
            w90=> c1_n0_w90, 
            w91=> c1_n0_w91, 
            w92=> c1_n0_w92, 
            w93=> c1_n0_w93, 
            w94=> c1_n0_w94, 
            w95=> c1_n0_w95, 
            w96=> c1_n0_w96, 
            w97=> c1_n0_w97, 
            w98=> c1_n0_w98, 
            w99=> c1_n0_w99, 
            w100=> c1_n0_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n0_y
   );           
            
neuron_inst_1: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n1_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n1_w1, 
            w2=> c1_n1_w2, 
            w3=> c1_n1_w3, 
            w4=> c1_n1_w4, 
            w5=> c1_n1_w5, 
            w6=> c1_n1_w6, 
            w7=> c1_n1_w7, 
            w8=> c1_n1_w8, 
            w9=> c1_n1_w9, 
            w10=> c1_n1_w10, 
            w11=> c1_n1_w11, 
            w12=> c1_n1_w12, 
            w13=> c1_n1_w13, 
            w14=> c1_n1_w14, 
            w15=> c1_n1_w15, 
            w16=> c1_n1_w16, 
            w17=> c1_n1_w17, 
            w18=> c1_n1_w18, 
            w19=> c1_n1_w19, 
            w20=> c1_n1_w20, 
            w21=> c1_n1_w21, 
            w22=> c1_n1_w22, 
            w23=> c1_n1_w23, 
            w24=> c1_n1_w24, 
            w25=> c1_n1_w25, 
            w26=> c1_n1_w26, 
            w27=> c1_n1_w27, 
            w28=> c1_n1_w28, 
            w29=> c1_n1_w29, 
            w30=> c1_n1_w30, 
            w31=> c1_n1_w31, 
            w32=> c1_n1_w32, 
            w33=> c1_n1_w33, 
            w34=> c1_n1_w34, 
            w35=> c1_n1_w35, 
            w36=> c1_n1_w36, 
            w37=> c1_n1_w37, 
            w38=> c1_n1_w38, 
            w39=> c1_n1_w39, 
            w40=> c1_n1_w40, 
            w41=> c1_n1_w41, 
            w42=> c1_n1_w42, 
            w43=> c1_n1_w43, 
            w44=> c1_n1_w44, 
            w45=> c1_n1_w45, 
            w46=> c1_n1_w46, 
            w47=> c1_n1_w47, 
            w48=> c1_n1_w48, 
            w49=> c1_n1_w49, 
            w50=> c1_n1_w50, 
            w51=> c1_n1_w51, 
            w52=> c1_n1_w52, 
            w53=> c1_n1_w53, 
            w54=> c1_n1_w54, 
            w55=> c1_n1_w55, 
            w56=> c1_n1_w56, 
            w57=> c1_n1_w57, 
            w58=> c1_n1_w58, 
            w59=> c1_n1_w59, 
            w60=> c1_n1_w60, 
            w61=> c1_n1_w61, 
            w62=> c1_n1_w62, 
            w63=> c1_n1_w63, 
            w64=> c1_n1_w64, 
            w65=> c1_n1_w65, 
            w66=> c1_n1_w66, 
            w67=> c1_n1_w67, 
            w68=> c1_n1_w68, 
            w69=> c1_n1_w69, 
            w70=> c1_n1_w70, 
            w71=> c1_n1_w71, 
            w72=> c1_n1_w72, 
            w73=> c1_n1_w73, 
            w74=> c1_n1_w74, 
            w75=> c1_n1_w75, 
            w76=> c1_n1_w76, 
            w77=> c1_n1_w77, 
            w78=> c1_n1_w78, 
            w79=> c1_n1_w79, 
            w80=> c1_n1_w80, 
            w81=> c1_n1_w81, 
            w82=> c1_n1_w82, 
            w83=> c1_n1_w83, 
            w84=> c1_n1_w84, 
            w85=> c1_n1_w85, 
            w86=> c1_n1_w86, 
            w87=> c1_n1_w87, 
            w88=> c1_n1_w88, 
            w89=> c1_n1_w89, 
            w90=> c1_n1_w90, 
            w91=> c1_n1_w91, 
            w92=> c1_n1_w92, 
            w93=> c1_n1_w93, 
            w94=> c1_n1_w94, 
            w95=> c1_n1_w95, 
            w96=> c1_n1_w96, 
            w97=> c1_n1_w97, 
            w98=> c1_n1_w98, 
            w99=> c1_n1_w99, 
            w100=> c1_n1_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n1_y
   );           
            
neuron_inst_2: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n2_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n2_w1, 
            w2=> c1_n2_w2, 
            w3=> c1_n2_w3, 
            w4=> c1_n2_w4, 
            w5=> c1_n2_w5, 
            w6=> c1_n2_w6, 
            w7=> c1_n2_w7, 
            w8=> c1_n2_w8, 
            w9=> c1_n2_w9, 
            w10=> c1_n2_w10, 
            w11=> c1_n2_w11, 
            w12=> c1_n2_w12, 
            w13=> c1_n2_w13, 
            w14=> c1_n2_w14, 
            w15=> c1_n2_w15, 
            w16=> c1_n2_w16, 
            w17=> c1_n2_w17, 
            w18=> c1_n2_w18, 
            w19=> c1_n2_w19, 
            w20=> c1_n2_w20, 
            w21=> c1_n2_w21, 
            w22=> c1_n2_w22, 
            w23=> c1_n2_w23, 
            w24=> c1_n2_w24, 
            w25=> c1_n2_w25, 
            w26=> c1_n2_w26, 
            w27=> c1_n2_w27, 
            w28=> c1_n2_w28, 
            w29=> c1_n2_w29, 
            w30=> c1_n2_w30, 
            w31=> c1_n2_w31, 
            w32=> c1_n2_w32, 
            w33=> c1_n2_w33, 
            w34=> c1_n2_w34, 
            w35=> c1_n2_w35, 
            w36=> c1_n2_w36, 
            w37=> c1_n2_w37, 
            w38=> c1_n2_w38, 
            w39=> c1_n2_w39, 
            w40=> c1_n2_w40, 
            w41=> c1_n2_w41, 
            w42=> c1_n2_w42, 
            w43=> c1_n2_w43, 
            w44=> c1_n2_w44, 
            w45=> c1_n2_w45, 
            w46=> c1_n2_w46, 
            w47=> c1_n2_w47, 
            w48=> c1_n2_w48, 
            w49=> c1_n2_w49, 
            w50=> c1_n2_w50, 
            w51=> c1_n2_w51, 
            w52=> c1_n2_w52, 
            w53=> c1_n2_w53, 
            w54=> c1_n2_w54, 
            w55=> c1_n2_w55, 
            w56=> c1_n2_w56, 
            w57=> c1_n2_w57, 
            w58=> c1_n2_w58, 
            w59=> c1_n2_w59, 
            w60=> c1_n2_w60, 
            w61=> c1_n2_w61, 
            w62=> c1_n2_w62, 
            w63=> c1_n2_w63, 
            w64=> c1_n2_w64, 
            w65=> c1_n2_w65, 
            w66=> c1_n2_w66, 
            w67=> c1_n2_w67, 
            w68=> c1_n2_w68, 
            w69=> c1_n2_w69, 
            w70=> c1_n2_w70, 
            w71=> c1_n2_w71, 
            w72=> c1_n2_w72, 
            w73=> c1_n2_w73, 
            w74=> c1_n2_w74, 
            w75=> c1_n2_w75, 
            w76=> c1_n2_w76, 
            w77=> c1_n2_w77, 
            w78=> c1_n2_w78, 
            w79=> c1_n2_w79, 
            w80=> c1_n2_w80, 
            w81=> c1_n2_w81, 
            w82=> c1_n2_w82, 
            w83=> c1_n2_w83, 
            w84=> c1_n2_w84, 
            w85=> c1_n2_w85, 
            w86=> c1_n2_w86, 
            w87=> c1_n2_w87, 
            w88=> c1_n2_w88, 
            w89=> c1_n2_w89, 
            w90=> c1_n2_w90, 
            w91=> c1_n2_w91, 
            w92=> c1_n2_w92, 
            w93=> c1_n2_w93, 
            w94=> c1_n2_w94, 
            w95=> c1_n2_w95, 
            w96=> c1_n2_w96, 
            w97=> c1_n2_w97, 
            w98=> c1_n2_w98, 
            w99=> c1_n2_w99, 
            w100=> c1_n2_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n2_y
   );           
            
neuron_inst_3: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n3_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n3_w1, 
            w2=> c1_n3_w2, 
            w3=> c1_n3_w3, 
            w4=> c1_n3_w4, 
            w5=> c1_n3_w5, 
            w6=> c1_n3_w6, 
            w7=> c1_n3_w7, 
            w8=> c1_n3_w8, 
            w9=> c1_n3_w9, 
            w10=> c1_n3_w10, 
            w11=> c1_n3_w11, 
            w12=> c1_n3_w12, 
            w13=> c1_n3_w13, 
            w14=> c1_n3_w14, 
            w15=> c1_n3_w15, 
            w16=> c1_n3_w16, 
            w17=> c1_n3_w17, 
            w18=> c1_n3_w18, 
            w19=> c1_n3_w19, 
            w20=> c1_n3_w20, 
            w21=> c1_n3_w21, 
            w22=> c1_n3_w22, 
            w23=> c1_n3_w23, 
            w24=> c1_n3_w24, 
            w25=> c1_n3_w25, 
            w26=> c1_n3_w26, 
            w27=> c1_n3_w27, 
            w28=> c1_n3_w28, 
            w29=> c1_n3_w29, 
            w30=> c1_n3_w30, 
            w31=> c1_n3_w31, 
            w32=> c1_n3_w32, 
            w33=> c1_n3_w33, 
            w34=> c1_n3_w34, 
            w35=> c1_n3_w35, 
            w36=> c1_n3_w36, 
            w37=> c1_n3_w37, 
            w38=> c1_n3_w38, 
            w39=> c1_n3_w39, 
            w40=> c1_n3_w40, 
            w41=> c1_n3_w41, 
            w42=> c1_n3_w42, 
            w43=> c1_n3_w43, 
            w44=> c1_n3_w44, 
            w45=> c1_n3_w45, 
            w46=> c1_n3_w46, 
            w47=> c1_n3_w47, 
            w48=> c1_n3_w48, 
            w49=> c1_n3_w49, 
            w50=> c1_n3_w50, 
            w51=> c1_n3_w51, 
            w52=> c1_n3_w52, 
            w53=> c1_n3_w53, 
            w54=> c1_n3_w54, 
            w55=> c1_n3_w55, 
            w56=> c1_n3_w56, 
            w57=> c1_n3_w57, 
            w58=> c1_n3_w58, 
            w59=> c1_n3_w59, 
            w60=> c1_n3_w60, 
            w61=> c1_n3_w61, 
            w62=> c1_n3_w62, 
            w63=> c1_n3_w63, 
            w64=> c1_n3_w64, 
            w65=> c1_n3_w65, 
            w66=> c1_n3_w66, 
            w67=> c1_n3_w67, 
            w68=> c1_n3_w68, 
            w69=> c1_n3_w69, 
            w70=> c1_n3_w70, 
            w71=> c1_n3_w71, 
            w72=> c1_n3_w72, 
            w73=> c1_n3_w73, 
            w74=> c1_n3_w74, 
            w75=> c1_n3_w75, 
            w76=> c1_n3_w76, 
            w77=> c1_n3_w77, 
            w78=> c1_n3_w78, 
            w79=> c1_n3_w79, 
            w80=> c1_n3_w80, 
            w81=> c1_n3_w81, 
            w82=> c1_n3_w82, 
            w83=> c1_n3_w83, 
            w84=> c1_n3_w84, 
            w85=> c1_n3_w85, 
            w86=> c1_n3_w86, 
            w87=> c1_n3_w87, 
            w88=> c1_n3_w88, 
            w89=> c1_n3_w89, 
            w90=> c1_n3_w90, 
            w91=> c1_n3_w91, 
            w92=> c1_n3_w92, 
            w93=> c1_n3_w93, 
            w94=> c1_n3_w94, 
            w95=> c1_n3_w95, 
            w96=> c1_n3_w96, 
            w97=> c1_n3_w97, 
            w98=> c1_n3_w98, 
            w99=> c1_n3_w99, 
            w100=> c1_n3_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n3_y
   );           
            
neuron_inst_4: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n4_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n4_w1, 
            w2=> c1_n4_w2, 
            w3=> c1_n4_w3, 
            w4=> c1_n4_w4, 
            w5=> c1_n4_w5, 
            w6=> c1_n4_w6, 
            w7=> c1_n4_w7, 
            w8=> c1_n4_w8, 
            w9=> c1_n4_w9, 
            w10=> c1_n4_w10, 
            w11=> c1_n4_w11, 
            w12=> c1_n4_w12, 
            w13=> c1_n4_w13, 
            w14=> c1_n4_w14, 
            w15=> c1_n4_w15, 
            w16=> c1_n4_w16, 
            w17=> c1_n4_w17, 
            w18=> c1_n4_w18, 
            w19=> c1_n4_w19, 
            w20=> c1_n4_w20, 
            w21=> c1_n4_w21, 
            w22=> c1_n4_w22, 
            w23=> c1_n4_w23, 
            w24=> c1_n4_w24, 
            w25=> c1_n4_w25, 
            w26=> c1_n4_w26, 
            w27=> c1_n4_w27, 
            w28=> c1_n4_w28, 
            w29=> c1_n4_w29, 
            w30=> c1_n4_w30, 
            w31=> c1_n4_w31, 
            w32=> c1_n4_w32, 
            w33=> c1_n4_w33, 
            w34=> c1_n4_w34, 
            w35=> c1_n4_w35, 
            w36=> c1_n4_w36, 
            w37=> c1_n4_w37, 
            w38=> c1_n4_w38, 
            w39=> c1_n4_w39, 
            w40=> c1_n4_w40, 
            w41=> c1_n4_w41, 
            w42=> c1_n4_w42, 
            w43=> c1_n4_w43, 
            w44=> c1_n4_w44, 
            w45=> c1_n4_w45, 
            w46=> c1_n4_w46, 
            w47=> c1_n4_w47, 
            w48=> c1_n4_w48, 
            w49=> c1_n4_w49, 
            w50=> c1_n4_w50, 
            w51=> c1_n4_w51, 
            w52=> c1_n4_w52, 
            w53=> c1_n4_w53, 
            w54=> c1_n4_w54, 
            w55=> c1_n4_w55, 
            w56=> c1_n4_w56, 
            w57=> c1_n4_w57, 
            w58=> c1_n4_w58, 
            w59=> c1_n4_w59, 
            w60=> c1_n4_w60, 
            w61=> c1_n4_w61, 
            w62=> c1_n4_w62, 
            w63=> c1_n4_w63, 
            w64=> c1_n4_w64, 
            w65=> c1_n4_w65, 
            w66=> c1_n4_w66, 
            w67=> c1_n4_w67, 
            w68=> c1_n4_w68, 
            w69=> c1_n4_w69, 
            w70=> c1_n4_w70, 
            w71=> c1_n4_w71, 
            w72=> c1_n4_w72, 
            w73=> c1_n4_w73, 
            w74=> c1_n4_w74, 
            w75=> c1_n4_w75, 
            w76=> c1_n4_w76, 
            w77=> c1_n4_w77, 
            w78=> c1_n4_w78, 
            w79=> c1_n4_w79, 
            w80=> c1_n4_w80, 
            w81=> c1_n4_w81, 
            w82=> c1_n4_w82, 
            w83=> c1_n4_w83, 
            w84=> c1_n4_w84, 
            w85=> c1_n4_w85, 
            w86=> c1_n4_w86, 
            w87=> c1_n4_w87, 
            w88=> c1_n4_w88, 
            w89=> c1_n4_w89, 
            w90=> c1_n4_w90, 
            w91=> c1_n4_w91, 
            w92=> c1_n4_w92, 
            w93=> c1_n4_w93, 
            w94=> c1_n4_w94, 
            w95=> c1_n4_w95, 
            w96=> c1_n4_w96, 
            w97=> c1_n4_w97, 
            w98=> c1_n4_w98, 
            w99=> c1_n4_w99, 
            w100=> c1_n4_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n4_y
   );           
            
neuron_inst_5: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n5_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n5_w1, 
            w2=> c1_n5_w2, 
            w3=> c1_n5_w3, 
            w4=> c1_n5_w4, 
            w5=> c1_n5_w5, 
            w6=> c1_n5_w6, 
            w7=> c1_n5_w7, 
            w8=> c1_n5_w8, 
            w9=> c1_n5_w9, 
            w10=> c1_n5_w10, 
            w11=> c1_n5_w11, 
            w12=> c1_n5_w12, 
            w13=> c1_n5_w13, 
            w14=> c1_n5_w14, 
            w15=> c1_n5_w15, 
            w16=> c1_n5_w16, 
            w17=> c1_n5_w17, 
            w18=> c1_n5_w18, 
            w19=> c1_n5_w19, 
            w20=> c1_n5_w20, 
            w21=> c1_n5_w21, 
            w22=> c1_n5_w22, 
            w23=> c1_n5_w23, 
            w24=> c1_n5_w24, 
            w25=> c1_n5_w25, 
            w26=> c1_n5_w26, 
            w27=> c1_n5_w27, 
            w28=> c1_n5_w28, 
            w29=> c1_n5_w29, 
            w30=> c1_n5_w30, 
            w31=> c1_n5_w31, 
            w32=> c1_n5_w32, 
            w33=> c1_n5_w33, 
            w34=> c1_n5_w34, 
            w35=> c1_n5_w35, 
            w36=> c1_n5_w36, 
            w37=> c1_n5_w37, 
            w38=> c1_n5_w38, 
            w39=> c1_n5_w39, 
            w40=> c1_n5_w40, 
            w41=> c1_n5_w41, 
            w42=> c1_n5_w42, 
            w43=> c1_n5_w43, 
            w44=> c1_n5_w44, 
            w45=> c1_n5_w45, 
            w46=> c1_n5_w46, 
            w47=> c1_n5_w47, 
            w48=> c1_n5_w48, 
            w49=> c1_n5_w49, 
            w50=> c1_n5_w50, 
            w51=> c1_n5_w51, 
            w52=> c1_n5_w52, 
            w53=> c1_n5_w53, 
            w54=> c1_n5_w54, 
            w55=> c1_n5_w55, 
            w56=> c1_n5_w56, 
            w57=> c1_n5_w57, 
            w58=> c1_n5_w58, 
            w59=> c1_n5_w59, 
            w60=> c1_n5_w60, 
            w61=> c1_n5_w61, 
            w62=> c1_n5_w62, 
            w63=> c1_n5_w63, 
            w64=> c1_n5_w64, 
            w65=> c1_n5_w65, 
            w66=> c1_n5_w66, 
            w67=> c1_n5_w67, 
            w68=> c1_n5_w68, 
            w69=> c1_n5_w69, 
            w70=> c1_n5_w70, 
            w71=> c1_n5_w71, 
            w72=> c1_n5_w72, 
            w73=> c1_n5_w73, 
            w74=> c1_n5_w74, 
            w75=> c1_n5_w75, 
            w76=> c1_n5_w76, 
            w77=> c1_n5_w77, 
            w78=> c1_n5_w78, 
            w79=> c1_n5_w79, 
            w80=> c1_n5_w80, 
            w81=> c1_n5_w81, 
            w82=> c1_n5_w82, 
            w83=> c1_n5_w83, 
            w84=> c1_n5_w84, 
            w85=> c1_n5_w85, 
            w86=> c1_n5_w86, 
            w87=> c1_n5_w87, 
            w88=> c1_n5_w88, 
            w89=> c1_n5_w89, 
            w90=> c1_n5_w90, 
            w91=> c1_n5_w91, 
            w92=> c1_n5_w92, 
            w93=> c1_n5_w93, 
            w94=> c1_n5_w94, 
            w95=> c1_n5_w95, 
            w96=> c1_n5_w96, 
            w97=> c1_n5_w97, 
            w98=> c1_n5_w98, 
            w99=> c1_n5_w99, 
            w100=> c1_n5_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n5_y
   );           
            
neuron_inst_6: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n6_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n6_w1, 
            w2=> c1_n6_w2, 
            w3=> c1_n6_w3, 
            w4=> c1_n6_w4, 
            w5=> c1_n6_w5, 
            w6=> c1_n6_w6, 
            w7=> c1_n6_w7, 
            w8=> c1_n6_w8, 
            w9=> c1_n6_w9, 
            w10=> c1_n6_w10, 
            w11=> c1_n6_w11, 
            w12=> c1_n6_w12, 
            w13=> c1_n6_w13, 
            w14=> c1_n6_w14, 
            w15=> c1_n6_w15, 
            w16=> c1_n6_w16, 
            w17=> c1_n6_w17, 
            w18=> c1_n6_w18, 
            w19=> c1_n6_w19, 
            w20=> c1_n6_w20, 
            w21=> c1_n6_w21, 
            w22=> c1_n6_w22, 
            w23=> c1_n6_w23, 
            w24=> c1_n6_w24, 
            w25=> c1_n6_w25, 
            w26=> c1_n6_w26, 
            w27=> c1_n6_w27, 
            w28=> c1_n6_w28, 
            w29=> c1_n6_w29, 
            w30=> c1_n6_w30, 
            w31=> c1_n6_w31, 
            w32=> c1_n6_w32, 
            w33=> c1_n6_w33, 
            w34=> c1_n6_w34, 
            w35=> c1_n6_w35, 
            w36=> c1_n6_w36, 
            w37=> c1_n6_w37, 
            w38=> c1_n6_w38, 
            w39=> c1_n6_w39, 
            w40=> c1_n6_w40, 
            w41=> c1_n6_w41, 
            w42=> c1_n6_w42, 
            w43=> c1_n6_w43, 
            w44=> c1_n6_w44, 
            w45=> c1_n6_w45, 
            w46=> c1_n6_w46, 
            w47=> c1_n6_w47, 
            w48=> c1_n6_w48, 
            w49=> c1_n6_w49, 
            w50=> c1_n6_w50, 
            w51=> c1_n6_w51, 
            w52=> c1_n6_w52, 
            w53=> c1_n6_w53, 
            w54=> c1_n6_w54, 
            w55=> c1_n6_w55, 
            w56=> c1_n6_w56, 
            w57=> c1_n6_w57, 
            w58=> c1_n6_w58, 
            w59=> c1_n6_w59, 
            w60=> c1_n6_w60, 
            w61=> c1_n6_w61, 
            w62=> c1_n6_w62, 
            w63=> c1_n6_w63, 
            w64=> c1_n6_w64, 
            w65=> c1_n6_w65, 
            w66=> c1_n6_w66, 
            w67=> c1_n6_w67, 
            w68=> c1_n6_w68, 
            w69=> c1_n6_w69, 
            w70=> c1_n6_w70, 
            w71=> c1_n6_w71, 
            w72=> c1_n6_w72, 
            w73=> c1_n6_w73, 
            w74=> c1_n6_w74, 
            w75=> c1_n6_w75, 
            w76=> c1_n6_w76, 
            w77=> c1_n6_w77, 
            w78=> c1_n6_w78, 
            w79=> c1_n6_w79, 
            w80=> c1_n6_w80, 
            w81=> c1_n6_w81, 
            w82=> c1_n6_w82, 
            w83=> c1_n6_w83, 
            w84=> c1_n6_w84, 
            w85=> c1_n6_w85, 
            w86=> c1_n6_w86, 
            w87=> c1_n6_w87, 
            w88=> c1_n6_w88, 
            w89=> c1_n6_w89, 
            w90=> c1_n6_w90, 
            w91=> c1_n6_w91, 
            w92=> c1_n6_w92, 
            w93=> c1_n6_w93, 
            w94=> c1_n6_w94, 
            w95=> c1_n6_w95, 
            w96=> c1_n6_w96, 
            w97=> c1_n6_w97, 
            w98=> c1_n6_w98, 
            w99=> c1_n6_w99, 
            w100=> c1_n6_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n6_y
   );           
            
neuron_inst_7: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n7_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n7_w1, 
            w2=> c1_n7_w2, 
            w3=> c1_n7_w3, 
            w4=> c1_n7_w4, 
            w5=> c1_n7_w5, 
            w6=> c1_n7_w6, 
            w7=> c1_n7_w7, 
            w8=> c1_n7_w8, 
            w9=> c1_n7_w9, 
            w10=> c1_n7_w10, 
            w11=> c1_n7_w11, 
            w12=> c1_n7_w12, 
            w13=> c1_n7_w13, 
            w14=> c1_n7_w14, 
            w15=> c1_n7_w15, 
            w16=> c1_n7_w16, 
            w17=> c1_n7_w17, 
            w18=> c1_n7_w18, 
            w19=> c1_n7_w19, 
            w20=> c1_n7_w20, 
            w21=> c1_n7_w21, 
            w22=> c1_n7_w22, 
            w23=> c1_n7_w23, 
            w24=> c1_n7_w24, 
            w25=> c1_n7_w25, 
            w26=> c1_n7_w26, 
            w27=> c1_n7_w27, 
            w28=> c1_n7_w28, 
            w29=> c1_n7_w29, 
            w30=> c1_n7_w30, 
            w31=> c1_n7_w31, 
            w32=> c1_n7_w32, 
            w33=> c1_n7_w33, 
            w34=> c1_n7_w34, 
            w35=> c1_n7_w35, 
            w36=> c1_n7_w36, 
            w37=> c1_n7_w37, 
            w38=> c1_n7_w38, 
            w39=> c1_n7_w39, 
            w40=> c1_n7_w40, 
            w41=> c1_n7_w41, 
            w42=> c1_n7_w42, 
            w43=> c1_n7_w43, 
            w44=> c1_n7_w44, 
            w45=> c1_n7_w45, 
            w46=> c1_n7_w46, 
            w47=> c1_n7_w47, 
            w48=> c1_n7_w48, 
            w49=> c1_n7_w49, 
            w50=> c1_n7_w50, 
            w51=> c1_n7_w51, 
            w52=> c1_n7_w52, 
            w53=> c1_n7_w53, 
            w54=> c1_n7_w54, 
            w55=> c1_n7_w55, 
            w56=> c1_n7_w56, 
            w57=> c1_n7_w57, 
            w58=> c1_n7_w58, 
            w59=> c1_n7_w59, 
            w60=> c1_n7_w60, 
            w61=> c1_n7_w61, 
            w62=> c1_n7_w62, 
            w63=> c1_n7_w63, 
            w64=> c1_n7_w64, 
            w65=> c1_n7_w65, 
            w66=> c1_n7_w66, 
            w67=> c1_n7_w67, 
            w68=> c1_n7_w68, 
            w69=> c1_n7_w69, 
            w70=> c1_n7_w70, 
            w71=> c1_n7_w71, 
            w72=> c1_n7_w72, 
            w73=> c1_n7_w73, 
            w74=> c1_n7_w74, 
            w75=> c1_n7_w75, 
            w76=> c1_n7_w76, 
            w77=> c1_n7_w77, 
            w78=> c1_n7_w78, 
            w79=> c1_n7_w79, 
            w80=> c1_n7_w80, 
            w81=> c1_n7_w81, 
            w82=> c1_n7_w82, 
            w83=> c1_n7_w83, 
            w84=> c1_n7_w84, 
            w85=> c1_n7_w85, 
            w86=> c1_n7_w86, 
            w87=> c1_n7_w87, 
            w88=> c1_n7_w88, 
            w89=> c1_n7_w89, 
            w90=> c1_n7_w90, 
            w91=> c1_n7_w91, 
            w92=> c1_n7_w92, 
            w93=> c1_n7_w93, 
            w94=> c1_n7_w94, 
            w95=> c1_n7_w95, 
            w96=> c1_n7_w96, 
            w97=> c1_n7_w97, 
            w98=> c1_n7_w98, 
            w99=> c1_n7_w99, 
            w100=> c1_n7_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n7_y
   );           
            
neuron_inst_8: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n8_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n8_w1, 
            w2=> c1_n8_w2, 
            w3=> c1_n8_w3, 
            w4=> c1_n8_w4, 
            w5=> c1_n8_w5, 
            w6=> c1_n8_w6, 
            w7=> c1_n8_w7, 
            w8=> c1_n8_w8, 
            w9=> c1_n8_w9, 
            w10=> c1_n8_w10, 
            w11=> c1_n8_w11, 
            w12=> c1_n8_w12, 
            w13=> c1_n8_w13, 
            w14=> c1_n8_w14, 
            w15=> c1_n8_w15, 
            w16=> c1_n8_w16, 
            w17=> c1_n8_w17, 
            w18=> c1_n8_w18, 
            w19=> c1_n8_w19, 
            w20=> c1_n8_w20, 
            w21=> c1_n8_w21, 
            w22=> c1_n8_w22, 
            w23=> c1_n8_w23, 
            w24=> c1_n8_w24, 
            w25=> c1_n8_w25, 
            w26=> c1_n8_w26, 
            w27=> c1_n8_w27, 
            w28=> c1_n8_w28, 
            w29=> c1_n8_w29, 
            w30=> c1_n8_w30, 
            w31=> c1_n8_w31, 
            w32=> c1_n8_w32, 
            w33=> c1_n8_w33, 
            w34=> c1_n8_w34, 
            w35=> c1_n8_w35, 
            w36=> c1_n8_w36, 
            w37=> c1_n8_w37, 
            w38=> c1_n8_w38, 
            w39=> c1_n8_w39, 
            w40=> c1_n8_w40, 
            w41=> c1_n8_w41, 
            w42=> c1_n8_w42, 
            w43=> c1_n8_w43, 
            w44=> c1_n8_w44, 
            w45=> c1_n8_w45, 
            w46=> c1_n8_w46, 
            w47=> c1_n8_w47, 
            w48=> c1_n8_w48, 
            w49=> c1_n8_w49, 
            w50=> c1_n8_w50, 
            w51=> c1_n8_w51, 
            w52=> c1_n8_w52, 
            w53=> c1_n8_w53, 
            w54=> c1_n8_w54, 
            w55=> c1_n8_w55, 
            w56=> c1_n8_w56, 
            w57=> c1_n8_w57, 
            w58=> c1_n8_w58, 
            w59=> c1_n8_w59, 
            w60=> c1_n8_w60, 
            w61=> c1_n8_w61, 
            w62=> c1_n8_w62, 
            w63=> c1_n8_w63, 
            w64=> c1_n8_w64, 
            w65=> c1_n8_w65, 
            w66=> c1_n8_w66, 
            w67=> c1_n8_w67, 
            w68=> c1_n8_w68, 
            w69=> c1_n8_w69, 
            w70=> c1_n8_w70, 
            w71=> c1_n8_w71, 
            w72=> c1_n8_w72, 
            w73=> c1_n8_w73, 
            w74=> c1_n8_w74, 
            w75=> c1_n8_w75, 
            w76=> c1_n8_w76, 
            w77=> c1_n8_w77, 
            w78=> c1_n8_w78, 
            w79=> c1_n8_w79, 
            w80=> c1_n8_w80, 
            w81=> c1_n8_w81, 
            w82=> c1_n8_w82, 
            w83=> c1_n8_w83, 
            w84=> c1_n8_w84, 
            w85=> c1_n8_w85, 
            w86=> c1_n8_w86, 
            w87=> c1_n8_w87, 
            w88=> c1_n8_w88, 
            w89=> c1_n8_w89, 
            w90=> c1_n8_w90, 
            w91=> c1_n8_w91, 
            w92=> c1_n8_w92, 
            w93=> c1_n8_w93, 
            w94=> c1_n8_w94, 
            w95=> c1_n8_w95, 
            w96=> c1_n8_w96, 
            w97=> c1_n8_w97, 
            w98=> c1_n8_w98, 
            w99=> c1_n8_w99, 
            w100=> c1_n8_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n8_y
   );           
            
neuron_inst_9: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n9_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n9_w1, 
            w2=> c1_n9_w2, 
            w3=> c1_n9_w3, 
            w4=> c1_n9_w4, 
            w5=> c1_n9_w5, 
            w6=> c1_n9_w6, 
            w7=> c1_n9_w7, 
            w8=> c1_n9_w8, 
            w9=> c1_n9_w9, 
            w10=> c1_n9_w10, 
            w11=> c1_n9_w11, 
            w12=> c1_n9_w12, 
            w13=> c1_n9_w13, 
            w14=> c1_n9_w14, 
            w15=> c1_n9_w15, 
            w16=> c1_n9_w16, 
            w17=> c1_n9_w17, 
            w18=> c1_n9_w18, 
            w19=> c1_n9_w19, 
            w20=> c1_n9_w20, 
            w21=> c1_n9_w21, 
            w22=> c1_n9_w22, 
            w23=> c1_n9_w23, 
            w24=> c1_n9_w24, 
            w25=> c1_n9_w25, 
            w26=> c1_n9_w26, 
            w27=> c1_n9_w27, 
            w28=> c1_n9_w28, 
            w29=> c1_n9_w29, 
            w30=> c1_n9_w30, 
            w31=> c1_n9_w31, 
            w32=> c1_n9_w32, 
            w33=> c1_n9_w33, 
            w34=> c1_n9_w34, 
            w35=> c1_n9_w35, 
            w36=> c1_n9_w36, 
            w37=> c1_n9_w37, 
            w38=> c1_n9_w38, 
            w39=> c1_n9_w39, 
            w40=> c1_n9_w40, 
            w41=> c1_n9_w41, 
            w42=> c1_n9_w42, 
            w43=> c1_n9_w43, 
            w44=> c1_n9_w44, 
            w45=> c1_n9_w45, 
            w46=> c1_n9_w46, 
            w47=> c1_n9_w47, 
            w48=> c1_n9_w48, 
            w49=> c1_n9_w49, 
            w50=> c1_n9_w50, 
            w51=> c1_n9_w51, 
            w52=> c1_n9_w52, 
            w53=> c1_n9_w53, 
            w54=> c1_n9_w54, 
            w55=> c1_n9_w55, 
            w56=> c1_n9_w56, 
            w57=> c1_n9_w57, 
            w58=> c1_n9_w58, 
            w59=> c1_n9_w59, 
            w60=> c1_n9_w60, 
            w61=> c1_n9_w61, 
            w62=> c1_n9_w62, 
            w63=> c1_n9_w63, 
            w64=> c1_n9_w64, 
            w65=> c1_n9_w65, 
            w66=> c1_n9_w66, 
            w67=> c1_n9_w67, 
            w68=> c1_n9_w68, 
            w69=> c1_n9_w69, 
            w70=> c1_n9_w70, 
            w71=> c1_n9_w71, 
            w72=> c1_n9_w72, 
            w73=> c1_n9_w73, 
            w74=> c1_n9_w74, 
            w75=> c1_n9_w75, 
            w76=> c1_n9_w76, 
            w77=> c1_n9_w77, 
            w78=> c1_n9_w78, 
            w79=> c1_n9_w79, 
            w80=> c1_n9_w80, 
            w81=> c1_n9_w81, 
            w82=> c1_n9_w82, 
            w83=> c1_n9_w83, 
            w84=> c1_n9_w84, 
            w85=> c1_n9_w85, 
            w86=> c1_n9_w86, 
            w87=> c1_n9_w87, 
            w88=> c1_n9_w88, 
            w89=> c1_n9_w89, 
            w90=> c1_n9_w90, 
            w91=> c1_n9_w91, 
            w92=> c1_n9_w92, 
            w93=> c1_n9_w93, 
            w94=> c1_n9_w94, 
            w95=> c1_n9_w95, 
            w96=> c1_n9_w96, 
            w97=> c1_n9_w97, 
            w98=> c1_n9_w98, 
            w99=> c1_n9_w99, 
            w100=> c1_n9_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n9_y
   );           
            
neuron_inst_10: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n10_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n10_w1, 
            w2=> c1_n10_w2, 
            w3=> c1_n10_w3, 
            w4=> c1_n10_w4, 
            w5=> c1_n10_w5, 
            w6=> c1_n10_w6, 
            w7=> c1_n10_w7, 
            w8=> c1_n10_w8, 
            w9=> c1_n10_w9, 
            w10=> c1_n10_w10, 
            w11=> c1_n10_w11, 
            w12=> c1_n10_w12, 
            w13=> c1_n10_w13, 
            w14=> c1_n10_w14, 
            w15=> c1_n10_w15, 
            w16=> c1_n10_w16, 
            w17=> c1_n10_w17, 
            w18=> c1_n10_w18, 
            w19=> c1_n10_w19, 
            w20=> c1_n10_w20, 
            w21=> c1_n10_w21, 
            w22=> c1_n10_w22, 
            w23=> c1_n10_w23, 
            w24=> c1_n10_w24, 
            w25=> c1_n10_w25, 
            w26=> c1_n10_w26, 
            w27=> c1_n10_w27, 
            w28=> c1_n10_w28, 
            w29=> c1_n10_w29, 
            w30=> c1_n10_w30, 
            w31=> c1_n10_w31, 
            w32=> c1_n10_w32, 
            w33=> c1_n10_w33, 
            w34=> c1_n10_w34, 
            w35=> c1_n10_w35, 
            w36=> c1_n10_w36, 
            w37=> c1_n10_w37, 
            w38=> c1_n10_w38, 
            w39=> c1_n10_w39, 
            w40=> c1_n10_w40, 
            w41=> c1_n10_w41, 
            w42=> c1_n10_w42, 
            w43=> c1_n10_w43, 
            w44=> c1_n10_w44, 
            w45=> c1_n10_w45, 
            w46=> c1_n10_w46, 
            w47=> c1_n10_w47, 
            w48=> c1_n10_w48, 
            w49=> c1_n10_w49, 
            w50=> c1_n10_w50, 
            w51=> c1_n10_w51, 
            w52=> c1_n10_w52, 
            w53=> c1_n10_w53, 
            w54=> c1_n10_w54, 
            w55=> c1_n10_w55, 
            w56=> c1_n10_w56, 
            w57=> c1_n10_w57, 
            w58=> c1_n10_w58, 
            w59=> c1_n10_w59, 
            w60=> c1_n10_w60, 
            w61=> c1_n10_w61, 
            w62=> c1_n10_w62, 
            w63=> c1_n10_w63, 
            w64=> c1_n10_w64, 
            w65=> c1_n10_w65, 
            w66=> c1_n10_w66, 
            w67=> c1_n10_w67, 
            w68=> c1_n10_w68, 
            w69=> c1_n10_w69, 
            w70=> c1_n10_w70, 
            w71=> c1_n10_w71, 
            w72=> c1_n10_w72, 
            w73=> c1_n10_w73, 
            w74=> c1_n10_w74, 
            w75=> c1_n10_w75, 
            w76=> c1_n10_w76, 
            w77=> c1_n10_w77, 
            w78=> c1_n10_w78, 
            w79=> c1_n10_w79, 
            w80=> c1_n10_w80, 
            w81=> c1_n10_w81, 
            w82=> c1_n10_w82, 
            w83=> c1_n10_w83, 
            w84=> c1_n10_w84, 
            w85=> c1_n10_w85, 
            w86=> c1_n10_w86, 
            w87=> c1_n10_w87, 
            w88=> c1_n10_w88, 
            w89=> c1_n10_w89, 
            w90=> c1_n10_w90, 
            w91=> c1_n10_w91, 
            w92=> c1_n10_w92, 
            w93=> c1_n10_w93, 
            w94=> c1_n10_w94, 
            w95=> c1_n10_w95, 
            w96=> c1_n10_w96, 
            w97=> c1_n10_w97, 
            w98=> c1_n10_w98, 
            w99=> c1_n10_w99, 
            w100=> c1_n10_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n10_y
   );           
            
neuron_inst_11: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n11_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n11_w1, 
            w2=> c1_n11_w2, 
            w3=> c1_n11_w3, 
            w4=> c1_n11_w4, 
            w5=> c1_n11_w5, 
            w6=> c1_n11_w6, 
            w7=> c1_n11_w7, 
            w8=> c1_n11_w8, 
            w9=> c1_n11_w9, 
            w10=> c1_n11_w10, 
            w11=> c1_n11_w11, 
            w12=> c1_n11_w12, 
            w13=> c1_n11_w13, 
            w14=> c1_n11_w14, 
            w15=> c1_n11_w15, 
            w16=> c1_n11_w16, 
            w17=> c1_n11_w17, 
            w18=> c1_n11_w18, 
            w19=> c1_n11_w19, 
            w20=> c1_n11_w20, 
            w21=> c1_n11_w21, 
            w22=> c1_n11_w22, 
            w23=> c1_n11_w23, 
            w24=> c1_n11_w24, 
            w25=> c1_n11_w25, 
            w26=> c1_n11_w26, 
            w27=> c1_n11_w27, 
            w28=> c1_n11_w28, 
            w29=> c1_n11_w29, 
            w30=> c1_n11_w30, 
            w31=> c1_n11_w31, 
            w32=> c1_n11_w32, 
            w33=> c1_n11_w33, 
            w34=> c1_n11_w34, 
            w35=> c1_n11_w35, 
            w36=> c1_n11_w36, 
            w37=> c1_n11_w37, 
            w38=> c1_n11_w38, 
            w39=> c1_n11_w39, 
            w40=> c1_n11_w40, 
            w41=> c1_n11_w41, 
            w42=> c1_n11_w42, 
            w43=> c1_n11_w43, 
            w44=> c1_n11_w44, 
            w45=> c1_n11_w45, 
            w46=> c1_n11_w46, 
            w47=> c1_n11_w47, 
            w48=> c1_n11_w48, 
            w49=> c1_n11_w49, 
            w50=> c1_n11_w50, 
            w51=> c1_n11_w51, 
            w52=> c1_n11_w52, 
            w53=> c1_n11_w53, 
            w54=> c1_n11_w54, 
            w55=> c1_n11_w55, 
            w56=> c1_n11_w56, 
            w57=> c1_n11_w57, 
            w58=> c1_n11_w58, 
            w59=> c1_n11_w59, 
            w60=> c1_n11_w60, 
            w61=> c1_n11_w61, 
            w62=> c1_n11_w62, 
            w63=> c1_n11_w63, 
            w64=> c1_n11_w64, 
            w65=> c1_n11_w65, 
            w66=> c1_n11_w66, 
            w67=> c1_n11_w67, 
            w68=> c1_n11_w68, 
            w69=> c1_n11_w69, 
            w70=> c1_n11_w70, 
            w71=> c1_n11_w71, 
            w72=> c1_n11_w72, 
            w73=> c1_n11_w73, 
            w74=> c1_n11_w74, 
            w75=> c1_n11_w75, 
            w76=> c1_n11_w76, 
            w77=> c1_n11_w77, 
            w78=> c1_n11_w78, 
            w79=> c1_n11_w79, 
            w80=> c1_n11_w80, 
            w81=> c1_n11_w81, 
            w82=> c1_n11_w82, 
            w83=> c1_n11_w83, 
            w84=> c1_n11_w84, 
            w85=> c1_n11_w85, 
            w86=> c1_n11_w86, 
            w87=> c1_n11_w87, 
            w88=> c1_n11_w88, 
            w89=> c1_n11_w89, 
            w90=> c1_n11_w90, 
            w91=> c1_n11_w91, 
            w92=> c1_n11_w92, 
            w93=> c1_n11_w93, 
            w94=> c1_n11_w94, 
            w95=> c1_n11_w95, 
            w96=> c1_n11_w96, 
            w97=> c1_n11_w97, 
            w98=> c1_n11_w98, 
            w99=> c1_n11_w99, 
            w100=> c1_n11_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n11_y
   );           
            
neuron_inst_12: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n12_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n12_w1, 
            w2=> c1_n12_w2, 
            w3=> c1_n12_w3, 
            w4=> c1_n12_w4, 
            w5=> c1_n12_w5, 
            w6=> c1_n12_w6, 
            w7=> c1_n12_w7, 
            w8=> c1_n12_w8, 
            w9=> c1_n12_w9, 
            w10=> c1_n12_w10, 
            w11=> c1_n12_w11, 
            w12=> c1_n12_w12, 
            w13=> c1_n12_w13, 
            w14=> c1_n12_w14, 
            w15=> c1_n12_w15, 
            w16=> c1_n12_w16, 
            w17=> c1_n12_w17, 
            w18=> c1_n12_w18, 
            w19=> c1_n12_w19, 
            w20=> c1_n12_w20, 
            w21=> c1_n12_w21, 
            w22=> c1_n12_w22, 
            w23=> c1_n12_w23, 
            w24=> c1_n12_w24, 
            w25=> c1_n12_w25, 
            w26=> c1_n12_w26, 
            w27=> c1_n12_w27, 
            w28=> c1_n12_w28, 
            w29=> c1_n12_w29, 
            w30=> c1_n12_w30, 
            w31=> c1_n12_w31, 
            w32=> c1_n12_w32, 
            w33=> c1_n12_w33, 
            w34=> c1_n12_w34, 
            w35=> c1_n12_w35, 
            w36=> c1_n12_w36, 
            w37=> c1_n12_w37, 
            w38=> c1_n12_w38, 
            w39=> c1_n12_w39, 
            w40=> c1_n12_w40, 
            w41=> c1_n12_w41, 
            w42=> c1_n12_w42, 
            w43=> c1_n12_w43, 
            w44=> c1_n12_w44, 
            w45=> c1_n12_w45, 
            w46=> c1_n12_w46, 
            w47=> c1_n12_w47, 
            w48=> c1_n12_w48, 
            w49=> c1_n12_w49, 
            w50=> c1_n12_w50, 
            w51=> c1_n12_w51, 
            w52=> c1_n12_w52, 
            w53=> c1_n12_w53, 
            w54=> c1_n12_w54, 
            w55=> c1_n12_w55, 
            w56=> c1_n12_w56, 
            w57=> c1_n12_w57, 
            w58=> c1_n12_w58, 
            w59=> c1_n12_w59, 
            w60=> c1_n12_w60, 
            w61=> c1_n12_w61, 
            w62=> c1_n12_w62, 
            w63=> c1_n12_w63, 
            w64=> c1_n12_w64, 
            w65=> c1_n12_w65, 
            w66=> c1_n12_w66, 
            w67=> c1_n12_w67, 
            w68=> c1_n12_w68, 
            w69=> c1_n12_w69, 
            w70=> c1_n12_w70, 
            w71=> c1_n12_w71, 
            w72=> c1_n12_w72, 
            w73=> c1_n12_w73, 
            w74=> c1_n12_w74, 
            w75=> c1_n12_w75, 
            w76=> c1_n12_w76, 
            w77=> c1_n12_w77, 
            w78=> c1_n12_w78, 
            w79=> c1_n12_w79, 
            w80=> c1_n12_w80, 
            w81=> c1_n12_w81, 
            w82=> c1_n12_w82, 
            w83=> c1_n12_w83, 
            w84=> c1_n12_w84, 
            w85=> c1_n12_w85, 
            w86=> c1_n12_w86, 
            w87=> c1_n12_w87, 
            w88=> c1_n12_w88, 
            w89=> c1_n12_w89, 
            w90=> c1_n12_w90, 
            w91=> c1_n12_w91, 
            w92=> c1_n12_w92, 
            w93=> c1_n12_w93, 
            w94=> c1_n12_w94, 
            w95=> c1_n12_w95, 
            w96=> c1_n12_w96, 
            w97=> c1_n12_w97, 
            w98=> c1_n12_w98, 
            w99=> c1_n12_w99, 
            w100=> c1_n12_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n12_y
   );           
            
neuron_inst_13: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n13_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n13_w1, 
            w2=> c1_n13_w2, 
            w3=> c1_n13_w3, 
            w4=> c1_n13_w4, 
            w5=> c1_n13_w5, 
            w6=> c1_n13_w6, 
            w7=> c1_n13_w7, 
            w8=> c1_n13_w8, 
            w9=> c1_n13_w9, 
            w10=> c1_n13_w10, 
            w11=> c1_n13_w11, 
            w12=> c1_n13_w12, 
            w13=> c1_n13_w13, 
            w14=> c1_n13_w14, 
            w15=> c1_n13_w15, 
            w16=> c1_n13_w16, 
            w17=> c1_n13_w17, 
            w18=> c1_n13_w18, 
            w19=> c1_n13_w19, 
            w20=> c1_n13_w20, 
            w21=> c1_n13_w21, 
            w22=> c1_n13_w22, 
            w23=> c1_n13_w23, 
            w24=> c1_n13_w24, 
            w25=> c1_n13_w25, 
            w26=> c1_n13_w26, 
            w27=> c1_n13_w27, 
            w28=> c1_n13_w28, 
            w29=> c1_n13_w29, 
            w30=> c1_n13_w30, 
            w31=> c1_n13_w31, 
            w32=> c1_n13_w32, 
            w33=> c1_n13_w33, 
            w34=> c1_n13_w34, 
            w35=> c1_n13_w35, 
            w36=> c1_n13_w36, 
            w37=> c1_n13_w37, 
            w38=> c1_n13_w38, 
            w39=> c1_n13_w39, 
            w40=> c1_n13_w40, 
            w41=> c1_n13_w41, 
            w42=> c1_n13_w42, 
            w43=> c1_n13_w43, 
            w44=> c1_n13_w44, 
            w45=> c1_n13_w45, 
            w46=> c1_n13_w46, 
            w47=> c1_n13_w47, 
            w48=> c1_n13_w48, 
            w49=> c1_n13_w49, 
            w50=> c1_n13_w50, 
            w51=> c1_n13_w51, 
            w52=> c1_n13_w52, 
            w53=> c1_n13_w53, 
            w54=> c1_n13_w54, 
            w55=> c1_n13_w55, 
            w56=> c1_n13_w56, 
            w57=> c1_n13_w57, 
            w58=> c1_n13_w58, 
            w59=> c1_n13_w59, 
            w60=> c1_n13_w60, 
            w61=> c1_n13_w61, 
            w62=> c1_n13_w62, 
            w63=> c1_n13_w63, 
            w64=> c1_n13_w64, 
            w65=> c1_n13_w65, 
            w66=> c1_n13_w66, 
            w67=> c1_n13_w67, 
            w68=> c1_n13_w68, 
            w69=> c1_n13_w69, 
            w70=> c1_n13_w70, 
            w71=> c1_n13_w71, 
            w72=> c1_n13_w72, 
            w73=> c1_n13_w73, 
            w74=> c1_n13_w74, 
            w75=> c1_n13_w75, 
            w76=> c1_n13_w76, 
            w77=> c1_n13_w77, 
            w78=> c1_n13_w78, 
            w79=> c1_n13_w79, 
            w80=> c1_n13_w80, 
            w81=> c1_n13_w81, 
            w82=> c1_n13_w82, 
            w83=> c1_n13_w83, 
            w84=> c1_n13_w84, 
            w85=> c1_n13_w85, 
            w86=> c1_n13_w86, 
            w87=> c1_n13_w87, 
            w88=> c1_n13_w88, 
            w89=> c1_n13_w89, 
            w90=> c1_n13_w90, 
            w91=> c1_n13_w91, 
            w92=> c1_n13_w92, 
            w93=> c1_n13_w93, 
            w94=> c1_n13_w94, 
            w95=> c1_n13_w95, 
            w96=> c1_n13_w96, 
            w97=> c1_n13_w97, 
            w98=> c1_n13_w98, 
            w99=> c1_n13_w99, 
            w100=> c1_n13_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n13_y
   );           
            
neuron_inst_14: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n14_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n14_w1, 
            w2=> c1_n14_w2, 
            w3=> c1_n14_w3, 
            w4=> c1_n14_w4, 
            w5=> c1_n14_w5, 
            w6=> c1_n14_w6, 
            w7=> c1_n14_w7, 
            w8=> c1_n14_w8, 
            w9=> c1_n14_w9, 
            w10=> c1_n14_w10, 
            w11=> c1_n14_w11, 
            w12=> c1_n14_w12, 
            w13=> c1_n14_w13, 
            w14=> c1_n14_w14, 
            w15=> c1_n14_w15, 
            w16=> c1_n14_w16, 
            w17=> c1_n14_w17, 
            w18=> c1_n14_w18, 
            w19=> c1_n14_w19, 
            w20=> c1_n14_w20, 
            w21=> c1_n14_w21, 
            w22=> c1_n14_w22, 
            w23=> c1_n14_w23, 
            w24=> c1_n14_w24, 
            w25=> c1_n14_w25, 
            w26=> c1_n14_w26, 
            w27=> c1_n14_w27, 
            w28=> c1_n14_w28, 
            w29=> c1_n14_w29, 
            w30=> c1_n14_w30, 
            w31=> c1_n14_w31, 
            w32=> c1_n14_w32, 
            w33=> c1_n14_w33, 
            w34=> c1_n14_w34, 
            w35=> c1_n14_w35, 
            w36=> c1_n14_w36, 
            w37=> c1_n14_w37, 
            w38=> c1_n14_w38, 
            w39=> c1_n14_w39, 
            w40=> c1_n14_w40, 
            w41=> c1_n14_w41, 
            w42=> c1_n14_w42, 
            w43=> c1_n14_w43, 
            w44=> c1_n14_w44, 
            w45=> c1_n14_w45, 
            w46=> c1_n14_w46, 
            w47=> c1_n14_w47, 
            w48=> c1_n14_w48, 
            w49=> c1_n14_w49, 
            w50=> c1_n14_w50, 
            w51=> c1_n14_w51, 
            w52=> c1_n14_w52, 
            w53=> c1_n14_w53, 
            w54=> c1_n14_w54, 
            w55=> c1_n14_w55, 
            w56=> c1_n14_w56, 
            w57=> c1_n14_w57, 
            w58=> c1_n14_w58, 
            w59=> c1_n14_w59, 
            w60=> c1_n14_w60, 
            w61=> c1_n14_w61, 
            w62=> c1_n14_w62, 
            w63=> c1_n14_w63, 
            w64=> c1_n14_w64, 
            w65=> c1_n14_w65, 
            w66=> c1_n14_w66, 
            w67=> c1_n14_w67, 
            w68=> c1_n14_w68, 
            w69=> c1_n14_w69, 
            w70=> c1_n14_w70, 
            w71=> c1_n14_w71, 
            w72=> c1_n14_w72, 
            w73=> c1_n14_w73, 
            w74=> c1_n14_w74, 
            w75=> c1_n14_w75, 
            w76=> c1_n14_w76, 
            w77=> c1_n14_w77, 
            w78=> c1_n14_w78, 
            w79=> c1_n14_w79, 
            w80=> c1_n14_w80, 
            w81=> c1_n14_w81, 
            w82=> c1_n14_w82, 
            w83=> c1_n14_w83, 
            w84=> c1_n14_w84, 
            w85=> c1_n14_w85, 
            w86=> c1_n14_w86, 
            w87=> c1_n14_w87, 
            w88=> c1_n14_w88, 
            w89=> c1_n14_w89, 
            w90=> c1_n14_w90, 
            w91=> c1_n14_w91, 
            w92=> c1_n14_w92, 
            w93=> c1_n14_w93, 
            w94=> c1_n14_w94, 
            w95=> c1_n14_w95, 
            w96=> c1_n14_w96, 
            w97=> c1_n14_w97, 
            w98=> c1_n14_w98, 
            w99=> c1_n14_w99, 
            w100=> c1_n14_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n14_y
   );           
            
neuron_inst_15: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n15_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n15_w1, 
            w2=> c1_n15_w2, 
            w3=> c1_n15_w3, 
            w4=> c1_n15_w4, 
            w5=> c1_n15_w5, 
            w6=> c1_n15_w6, 
            w7=> c1_n15_w7, 
            w8=> c1_n15_w8, 
            w9=> c1_n15_w9, 
            w10=> c1_n15_w10, 
            w11=> c1_n15_w11, 
            w12=> c1_n15_w12, 
            w13=> c1_n15_w13, 
            w14=> c1_n15_w14, 
            w15=> c1_n15_w15, 
            w16=> c1_n15_w16, 
            w17=> c1_n15_w17, 
            w18=> c1_n15_w18, 
            w19=> c1_n15_w19, 
            w20=> c1_n15_w20, 
            w21=> c1_n15_w21, 
            w22=> c1_n15_w22, 
            w23=> c1_n15_w23, 
            w24=> c1_n15_w24, 
            w25=> c1_n15_w25, 
            w26=> c1_n15_w26, 
            w27=> c1_n15_w27, 
            w28=> c1_n15_w28, 
            w29=> c1_n15_w29, 
            w30=> c1_n15_w30, 
            w31=> c1_n15_w31, 
            w32=> c1_n15_w32, 
            w33=> c1_n15_w33, 
            w34=> c1_n15_w34, 
            w35=> c1_n15_w35, 
            w36=> c1_n15_w36, 
            w37=> c1_n15_w37, 
            w38=> c1_n15_w38, 
            w39=> c1_n15_w39, 
            w40=> c1_n15_w40, 
            w41=> c1_n15_w41, 
            w42=> c1_n15_w42, 
            w43=> c1_n15_w43, 
            w44=> c1_n15_w44, 
            w45=> c1_n15_w45, 
            w46=> c1_n15_w46, 
            w47=> c1_n15_w47, 
            w48=> c1_n15_w48, 
            w49=> c1_n15_w49, 
            w50=> c1_n15_w50, 
            w51=> c1_n15_w51, 
            w52=> c1_n15_w52, 
            w53=> c1_n15_w53, 
            w54=> c1_n15_w54, 
            w55=> c1_n15_w55, 
            w56=> c1_n15_w56, 
            w57=> c1_n15_w57, 
            w58=> c1_n15_w58, 
            w59=> c1_n15_w59, 
            w60=> c1_n15_w60, 
            w61=> c1_n15_w61, 
            w62=> c1_n15_w62, 
            w63=> c1_n15_w63, 
            w64=> c1_n15_w64, 
            w65=> c1_n15_w65, 
            w66=> c1_n15_w66, 
            w67=> c1_n15_w67, 
            w68=> c1_n15_w68, 
            w69=> c1_n15_w69, 
            w70=> c1_n15_w70, 
            w71=> c1_n15_w71, 
            w72=> c1_n15_w72, 
            w73=> c1_n15_w73, 
            w74=> c1_n15_w74, 
            w75=> c1_n15_w75, 
            w76=> c1_n15_w76, 
            w77=> c1_n15_w77, 
            w78=> c1_n15_w78, 
            w79=> c1_n15_w79, 
            w80=> c1_n15_w80, 
            w81=> c1_n15_w81, 
            w82=> c1_n15_w82, 
            w83=> c1_n15_w83, 
            w84=> c1_n15_w84, 
            w85=> c1_n15_w85, 
            w86=> c1_n15_w86, 
            w87=> c1_n15_w87, 
            w88=> c1_n15_w88, 
            w89=> c1_n15_w89, 
            w90=> c1_n15_w90, 
            w91=> c1_n15_w91, 
            w92=> c1_n15_w92, 
            w93=> c1_n15_w93, 
            w94=> c1_n15_w94, 
            w95=> c1_n15_w95, 
            w96=> c1_n15_w96, 
            w97=> c1_n15_w97, 
            w98=> c1_n15_w98, 
            w99=> c1_n15_w99, 
            w100=> c1_n15_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n15_y
   );           
            
neuron_inst_16: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n16_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n16_w1, 
            w2=> c1_n16_w2, 
            w3=> c1_n16_w3, 
            w4=> c1_n16_w4, 
            w5=> c1_n16_w5, 
            w6=> c1_n16_w6, 
            w7=> c1_n16_w7, 
            w8=> c1_n16_w8, 
            w9=> c1_n16_w9, 
            w10=> c1_n16_w10, 
            w11=> c1_n16_w11, 
            w12=> c1_n16_w12, 
            w13=> c1_n16_w13, 
            w14=> c1_n16_w14, 
            w15=> c1_n16_w15, 
            w16=> c1_n16_w16, 
            w17=> c1_n16_w17, 
            w18=> c1_n16_w18, 
            w19=> c1_n16_w19, 
            w20=> c1_n16_w20, 
            w21=> c1_n16_w21, 
            w22=> c1_n16_w22, 
            w23=> c1_n16_w23, 
            w24=> c1_n16_w24, 
            w25=> c1_n16_w25, 
            w26=> c1_n16_w26, 
            w27=> c1_n16_w27, 
            w28=> c1_n16_w28, 
            w29=> c1_n16_w29, 
            w30=> c1_n16_w30, 
            w31=> c1_n16_w31, 
            w32=> c1_n16_w32, 
            w33=> c1_n16_w33, 
            w34=> c1_n16_w34, 
            w35=> c1_n16_w35, 
            w36=> c1_n16_w36, 
            w37=> c1_n16_w37, 
            w38=> c1_n16_w38, 
            w39=> c1_n16_w39, 
            w40=> c1_n16_w40, 
            w41=> c1_n16_w41, 
            w42=> c1_n16_w42, 
            w43=> c1_n16_w43, 
            w44=> c1_n16_w44, 
            w45=> c1_n16_w45, 
            w46=> c1_n16_w46, 
            w47=> c1_n16_w47, 
            w48=> c1_n16_w48, 
            w49=> c1_n16_w49, 
            w50=> c1_n16_w50, 
            w51=> c1_n16_w51, 
            w52=> c1_n16_w52, 
            w53=> c1_n16_w53, 
            w54=> c1_n16_w54, 
            w55=> c1_n16_w55, 
            w56=> c1_n16_w56, 
            w57=> c1_n16_w57, 
            w58=> c1_n16_w58, 
            w59=> c1_n16_w59, 
            w60=> c1_n16_w60, 
            w61=> c1_n16_w61, 
            w62=> c1_n16_w62, 
            w63=> c1_n16_w63, 
            w64=> c1_n16_w64, 
            w65=> c1_n16_w65, 
            w66=> c1_n16_w66, 
            w67=> c1_n16_w67, 
            w68=> c1_n16_w68, 
            w69=> c1_n16_w69, 
            w70=> c1_n16_w70, 
            w71=> c1_n16_w71, 
            w72=> c1_n16_w72, 
            w73=> c1_n16_w73, 
            w74=> c1_n16_w74, 
            w75=> c1_n16_w75, 
            w76=> c1_n16_w76, 
            w77=> c1_n16_w77, 
            w78=> c1_n16_w78, 
            w79=> c1_n16_w79, 
            w80=> c1_n16_w80, 
            w81=> c1_n16_w81, 
            w82=> c1_n16_w82, 
            w83=> c1_n16_w83, 
            w84=> c1_n16_w84, 
            w85=> c1_n16_w85, 
            w86=> c1_n16_w86, 
            w87=> c1_n16_w87, 
            w88=> c1_n16_w88, 
            w89=> c1_n16_w89, 
            w90=> c1_n16_w90, 
            w91=> c1_n16_w91, 
            w92=> c1_n16_w92, 
            w93=> c1_n16_w93, 
            w94=> c1_n16_w94, 
            w95=> c1_n16_w95, 
            w96=> c1_n16_w96, 
            w97=> c1_n16_w97, 
            w98=> c1_n16_w98, 
            w99=> c1_n16_w99, 
            w100=> c1_n16_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n16_y
   );           
            
neuron_inst_17: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n17_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n17_w1, 
            w2=> c1_n17_w2, 
            w3=> c1_n17_w3, 
            w4=> c1_n17_w4, 
            w5=> c1_n17_w5, 
            w6=> c1_n17_w6, 
            w7=> c1_n17_w7, 
            w8=> c1_n17_w8, 
            w9=> c1_n17_w9, 
            w10=> c1_n17_w10, 
            w11=> c1_n17_w11, 
            w12=> c1_n17_w12, 
            w13=> c1_n17_w13, 
            w14=> c1_n17_w14, 
            w15=> c1_n17_w15, 
            w16=> c1_n17_w16, 
            w17=> c1_n17_w17, 
            w18=> c1_n17_w18, 
            w19=> c1_n17_w19, 
            w20=> c1_n17_w20, 
            w21=> c1_n17_w21, 
            w22=> c1_n17_w22, 
            w23=> c1_n17_w23, 
            w24=> c1_n17_w24, 
            w25=> c1_n17_w25, 
            w26=> c1_n17_w26, 
            w27=> c1_n17_w27, 
            w28=> c1_n17_w28, 
            w29=> c1_n17_w29, 
            w30=> c1_n17_w30, 
            w31=> c1_n17_w31, 
            w32=> c1_n17_w32, 
            w33=> c1_n17_w33, 
            w34=> c1_n17_w34, 
            w35=> c1_n17_w35, 
            w36=> c1_n17_w36, 
            w37=> c1_n17_w37, 
            w38=> c1_n17_w38, 
            w39=> c1_n17_w39, 
            w40=> c1_n17_w40, 
            w41=> c1_n17_w41, 
            w42=> c1_n17_w42, 
            w43=> c1_n17_w43, 
            w44=> c1_n17_w44, 
            w45=> c1_n17_w45, 
            w46=> c1_n17_w46, 
            w47=> c1_n17_w47, 
            w48=> c1_n17_w48, 
            w49=> c1_n17_w49, 
            w50=> c1_n17_w50, 
            w51=> c1_n17_w51, 
            w52=> c1_n17_w52, 
            w53=> c1_n17_w53, 
            w54=> c1_n17_w54, 
            w55=> c1_n17_w55, 
            w56=> c1_n17_w56, 
            w57=> c1_n17_w57, 
            w58=> c1_n17_w58, 
            w59=> c1_n17_w59, 
            w60=> c1_n17_w60, 
            w61=> c1_n17_w61, 
            w62=> c1_n17_w62, 
            w63=> c1_n17_w63, 
            w64=> c1_n17_w64, 
            w65=> c1_n17_w65, 
            w66=> c1_n17_w66, 
            w67=> c1_n17_w67, 
            w68=> c1_n17_w68, 
            w69=> c1_n17_w69, 
            w70=> c1_n17_w70, 
            w71=> c1_n17_w71, 
            w72=> c1_n17_w72, 
            w73=> c1_n17_w73, 
            w74=> c1_n17_w74, 
            w75=> c1_n17_w75, 
            w76=> c1_n17_w76, 
            w77=> c1_n17_w77, 
            w78=> c1_n17_w78, 
            w79=> c1_n17_w79, 
            w80=> c1_n17_w80, 
            w81=> c1_n17_w81, 
            w82=> c1_n17_w82, 
            w83=> c1_n17_w83, 
            w84=> c1_n17_w84, 
            w85=> c1_n17_w85, 
            w86=> c1_n17_w86, 
            w87=> c1_n17_w87, 
            w88=> c1_n17_w88, 
            w89=> c1_n17_w89, 
            w90=> c1_n17_w90, 
            w91=> c1_n17_w91, 
            w92=> c1_n17_w92, 
            w93=> c1_n17_w93, 
            w94=> c1_n17_w94, 
            w95=> c1_n17_w95, 
            w96=> c1_n17_w96, 
            w97=> c1_n17_w97, 
            w98=> c1_n17_w98, 
            w99=> c1_n17_w99, 
            w100=> c1_n17_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n17_y
   );           
            
neuron_inst_18: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n18_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n18_w1, 
            w2=> c1_n18_w2, 
            w3=> c1_n18_w3, 
            w4=> c1_n18_w4, 
            w5=> c1_n18_w5, 
            w6=> c1_n18_w6, 
            w7=> c1_n18_w7, 
            w8=> c1_n18_w8, 
            w9=> c1_n18_w9, 
            w10=> c1_n18_w10, 
            w11=> c1_n18_w11, 
            w12=> c1_n18_w12, 
            w13=> c1_n18_w13, 
            w14=> c1_n18_w14, 
            w15=> c1_n18_w15, 
            w16=> c1_n18_w16, 
            w17=> c1_n18_w17, 
            w18=> c1_n18_w18, 
            w19=> c1_n18_w19, 
            w20=> c1_n18_w20, 
            w21=> c1_n18_w21, 
            w22=> c1_n18_w22, 
            w23=> c1_n18_w23, 
            w24=> c1_n18_w24, 
            w25=> c1_n18_w25, 
            w26=> c1_n18_w26, 
            w27=> c1_n18_w27, 
            w28=> c1_n18_w28, 
            w29=> c1_n18_w29, 
            w30=> c1_n18_w30, 
            w31=> c1_n18_w31, 
            w32=> c1_n18_w32, 
            w33=> c1_n18_w33, 
            w34=> c1_n18_w34, 
            w35=> c1_n18_w35, 
            w36=> c1_n18_w36, 
            w37=> c1_n18_w37, 
            w38=> c1_n18_w38, 
            w39=> c1_n18_w39, 
            w40=> c1_n18_w40, 
            w41=> c1_n18_w41, 
            w42=> c1_n18_w42, 
            w43=> c1_n18_w43, 
            w44=> c1_n18_w44, 
            w45=> c1_n18_w45, 
            w46=> c1_n18_w46, 
            w47=> c1_n18_w47, 
            w48=> c1_n18_w48, 
            w49=> c1_n18_w49, 
            w50=> c1_n18_w50, 
            w51=> c1_n18_w51, 
            w52=> c1_n18_w52, 
            w53=> c1_n18_w53, 
            w54=> c1_n18_w54, 
            w55=> c1_n18_w55, 
            w56=> c1_n18_w56, 
            w57=> c1_n18_w57, 
            w58=> c1_n18_w58, 
            w59=> c1_n18_w59, 
            w60=> c1_n18_w60, 
            w61=> c1_n18_w61, 
            w62=> c1_n18_w62, 
            w63=> c1_n18_w63, 
            w64=> c1_n18_w64, 
            w65=> c1_n18_w65, 
            w66=> c1_n18_w66, 
            w67=> c1_n18_w67, 
            w68=> c1_n18_w68, 
            w69=> c1_n18_w69, 
            w70=> c1_n18_w70, 
            w71=> c1_n18_w71, 
            w72=> c1_n18_w72, 
            w73=> c1_n18_w73, 
            w74=> c1_n18_w74, 
            w75=> c1_n18_w75, 
            w76=> c1_n18_w76, 
            w77=> c1_n18_w77, 
            w78=> c1_n18_w78, 
            w79=> c1_n18_w79, 
            w80=> c1_n18_w80, 
            w81=> c1_n18_w81, 
            w82=> c1_n18_w82, 
            w83=> c1_n18_w83, 
            w84=> c1_n18_w84, 
            w85=> c1_n18_w85, 
            w86=> c1_n18_w86, 
            w87=> c1_n18_w87, 
            w88=> c1_n18_w88, 
            w89=> c1_n18_w89, 
            w90=> c1_n18_w90, 
            w91=> c1_n18_w91, 
            w92=> c1_n18_w92, 
            w93=> c1_n18_w93, 
            w94=> c1_n18_w94, 
            w95=> c1_n18_w95, 
            w96=> c1_n18_w96, 
            w97=> c1_n18_w97, 
            w98=> c1_n18_w98, 
            w99=> c1_n18_w99, 
            w100=> c1_n18_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n18_y
   );           
            
neuron_inst_19: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n19_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n19_w1, 
            w2=> c1_n19_w2, 
            w3=> c1_n19_w3, 
            w4=> c1_n19_w4, 
            w5=> c1_n19_w5, 
            w6=> c1_n19_w6, 
            w7=> c1_n19_w7, 
            w8=> c1_n19_w8, 
            w9=> c1_n19_w9, 
            w10=> c1_n19_w10, 
            w11=> c1_n19_w11, 
            w12=> c1_n19_w12, 
            w13=> c1_n19_w13, 
            w14=> c1_n19_w14, 
            w15=> c1_n19_w15, 
            w16=> c1_n19_w16, 
            w17=> c1_n19_w17, 
            w18=> c1_n19_w18, 
            w19=> c1_n19_w19, 
            w20=> c1_n19_w20, 
            w21=> c1_n19_w21, 
            w22=> c1_n19_w22, 
            w23=> c1_n19_w23, 
            w24=> c1_n19_w24, 
            w25=> c1_n19_w25, 
            w26=> c1_n19_w26, 
            w27=> c1_n19_w27, 
            w28=> c1_n19_w28, 
            w29=> c1_n19_w29, 
            w30=> c1_n19_w30, 
            w31=> c1_n19_w31, 
            w32=> c1_n19_w32, 
            w33=> c1_n19_w33, 
            w34=> c1_n19_w34, 
            w35=> c1_n19_w35, 
            w36=> c1_n19_w36, 
            w37=> c1_n19_w37, 
            w38=> c1_n19_w38, 
            w39=> c1_n19_w39, 
            w40=> c1_n19_w40, 
            w41=> c1_n19_w41, 
            w42=> c1_n19_w42, 
            w43=> c1_n19_w43, 
            w44=> c1_n19_w44, 
            w45=> c1_n19_w45, 
            w46=> c1_n19_w46, 
            w47=> c1_n19_w47, 
            w48=> c1_n19_w48, 
            w49=> c1_n19_w49, 
            w50=> c1_n19_w50, 
            w51=> c1_n19_w51, 
            w52=> c1_n19_w52, 
            w53=> c1_n19_w53, 
            w54=> c1_n19_w54, 
            w55=> c1_n19_w55, 
            w56=> c1_n19_w56, 
            w57=> c1_n19_w57, 
            w58=> c1_n19_w58, 
            w59=> c1_n19_w59, 
            w60=> c1_n19_w60, 
            w61=> c1_n19_w61, 
            w62=> c1_n19_w62, 
            w63=> c1_n19_w63, 
            w64=> c1_n19_w64, 
            w65=> c1_n19_w65, 
            w66=> c1_n19_w66, 
            w67=> c1_n19_w67, 
            w68=> c1_n19_w68, 
            w69=> c1_n19_w69, 
            w70=> c1_n19_w70, 
            w71=> c1_n19_w71, 
            w72=> c1_n19_w72, 
            w73=> c1_n19_w73, 
            w74=> c1_n19_w74, 
            w75=> c1_n19_w75, 
            w76=> c1_n19_w76, 
            w77=> c1_n19_w77, 
            w78=> c1_n19_w78, 
            w79=> c1_n19_w79, 
            w80=> c1_n19_w80, 
            w81=> c1_n19_w81, 
            w82=> c1_n19_w82, 
            w83=> c1_n19_w83, 
            w84=> c1_n19_w84, 
            w85=> c1_n19_w85, 
            w86=> c1_n19_w86, 
            w87=> c1_n19_w87, 
            w88=> c1_n19_w88, 
            w89=> c1_n19_w89, 
            w90=> c1_n19_w90, 
            w91=> c1_n19_w91, 
            w92=> c1_n19_w92, 
            w93=> c1_n19_w93, 
            w94=> c1_n19_w94, 
            w95=> c1_n19_w95, 
            w96=> c1_n19_w96, 
            w97=> c1_n19_w97, 
            w98=> c1_n19_w98, 
            w99=> c1_n19_w99, 
            w100=> c1_n19_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n19_y
   );           
            
neuron_inst_20: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n20_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n20_w1, 
            w2=> c1_n20_w2, 
            w3=> c1_n20_w3, 
            w4=> c1_n20_w4, 
            w5=> c1_n20_w5, 
            w6=> c1_n20_w6, 
            w7=> c1_n20_w7, 
            w8=> c1_n20_w8, 
            w9=> c1_n20_w9, 
            w10=> c1_n20_w10, 
            w11=> c1_n20_w11, 
            w12=> c1_n20_w12, 
            w13=> c1_n20_w13, 
            w14=> c1_n20_w14, 
            w15=> c1_n20_w15, 
            w16=> c1_n20_w16, 
            w17=> c1_n20_w17, 
            w18=> c1_n20_w18, 
            w19=> c1_n20_w19, 
            w20=> c1_n20_w20, 
            w21=> c1_n20_w21, 
            w22=> c1_n20_w22, 
            w23=> c1_n20_w23, 
            w24=> c1_n20_w24, 
            w25=> c1_n20_w25, 
            w26=> c1_n20_w26, 
            w27=> c1_n20_w27, 
            w28=> c1_n20_w28, 
            w29=> c1_n20_w29, 
            w30=> c1_n20_w30, 
            w31=> c1_n20_w31, 
            w32=> c1_n20_w32, 
            w33=> c1_n20_w33, 
            w34=> c1_n20_w34, 
            w35=> c1_n20_w35, 
            w36=> c1_n20_w36, 
            w37=> c1_n20_w37, 
            w38=> c1_n20_w38, 
            w39=> c1_n20_w39, 
            w40=> c1_n20_w40, 
            w41=> c1_n20_w41, 
            w42=> c1_n20_w42, 
            w43=> c1_n20_w43, 
            w44=> c1_n20_w44, 
            w45=> c1_n20_w45, 
            w46=> c1_n20_w46, 
            w47=> c1_n20_w47, 
            w48=> c1_n20_w48, 
            w49=> c1_n20_w49, 
            w50=> c1_n20_w50, 
            w51=> c1_n20_w51, 
            w52=> c1_n20_w52, 
            w53=> c1_n20_w53, 
            w54=> c1_n20_w54, 
            w55=> c1_n20_w55, 
            w56=> c1_n20_w56, 
            w57=> c1_n20_w57, 
            w58=> c1_n20_w58, 
            w59=> c1_n20_w59, 
            w60=> c1_n20_w60, 
            w61=> c1_n20_w61, 
            w62=> c1_n20_w62, 
            w63=> c1_n20_w63, 
            w64=> c1_n20_w64, 
            w65=> c1_n20_w65, 
            w66=> c1_n20_w66, 
            w67=> c1_n20_w67, 
            w68=> c1_n20_w68, 
            w69=> c1_n20_w69, 
            w70=> c1_n20_w70, 
            w71=> c1_n20_w71, 
            w72=> c1_n20_w72, 
            w73=> c1_n20_w73, 
            w74=> c1_n20_w74, 
            w75=> c1_n20_w75, 
            w76=> c1_n20_w76, 
            w77=> c1_n20_w77, 
            w78=> c1_n20_w78, 
            w79=> c1_n20_w79, 
            w80=> c1_n20_w80, 
            w81=> c1_n20_w81, 
            w82=> c1_n20_w82, 
            w83=> c1_n20_w83, 
            w84=> c1_n20_w84, 
            w85=> c1_n20_w85, 
            w86=> c1_n20_w86, 
            w87=> c1_n20_w87, 
            w88=> c1_n20_w88, 
            w89=> c1_n20_w89, 
            w90=> c1_n20_w90, 
            w91=> c1_n20_w91, 
            w92=> c1_n20_w92, 
            w93=> c1_n20_w93, 
            w94=> c1_n20_w94, 
            w95=> c1_n20_w95, 
            w96=> c1_n20_w96, 
            w97=> c1_n20_w97, 
            w98=> c1_n20_w98, 
            w99=> c1_n20_w99, 
            w100=> c1_n20_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n20_y
   );           
            
neuron_inst_21: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n21_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n21_w1, 
            w2=> c1_n21_w2, 
            w3=> c1_n21_w3, 
            w4=> c1_n21_w4, 
            w5=> c1_n21_w5, 
            w6=> c1_n21_w6, 
            w7=> c1_n21_w7, 
            w8=> c1_n21_w8, 
            w9=> c1_n21_w9, 
            w10=> c1_n21_w10, 
            w11=> c1_n21_w11, 
            w12=> c1_n21_w12, 
            w13=> c1_n21_w13, 
            w14=> c1_n21_w14, 
            w15=> c1_n21_w15, 
            w16=> c1_n21_w16, 
            w17=> c1_n21_w17, 
            w18=> c1_n21_w18, 
            w19=> c1_n21_w19, 
            w20=> c1_n21_w20, 
            w21=> c1_n21_w21, 
            w22=> c1_n21_w22, 
            w23=> c1_n21_w23, 
            w24=> c1_n21_w24, 
            w25=> c1_n21_w25, 
            w26=> c1_n21_w26, 
            w27=> c1_n21_w27, 
            w28=> c1_n21_w28, 
            w29=> c1_n21_w29, 
            w30=> c1_n21_w30, 
            w31=> c1_n21_w31, 
            w32=> c1_n21_w32, 
            w33=> c1_n21_w33, 
            w34=> c1_n21_w34, 
            w35=> c1_n21_w35, 
            w36=> c1_n21_w36, 
            w37=> c1_n21_w37, 
            w38=> c1_n21_w38, 
            w39=> c1_n21_w39, 
            w40=> c1_n21_w40, 
            w41=> c1_n21_w41, 
            w42=> c1_n21_w42, 
            w43=> c1_n21_w43, 
            w44=> c1_n21_w44, 
            w45=> c1_n21_w45, 
            w46=> c1_n21_w46, 
            w47=> c1_n21_w47, 
            w48=> c1_n21_w48, 
            w49=> c1_n21_w49, 
            w50=> c1_n21_w50, 
            w51=> c1_n21_w51, 
            w52=> c1_n21_w52, 
            w53=> c1_n21_w53, 
            w54=> c1_n21_w54, 
            w55=> c1_n21_w55, 
            w56=> c1_n21_w56, 
            w57=> c1_n21_w57, 
            w58=> c1_n21_w58, 
            w59=> c1_n21_w59, 
            w60=> c1_n21_w60, 
            w61=> c1_n21_w61, 
            w62=> c1_n21_w62, 
            w63=> c1_n21_w63, 
            w64=> c1_n21_w64, 
            w65=> c1_n21_w65, 
            w66=> c1_n21_w66, 
            w67=> c1_n21_w67, 
            w68=> c1_n21_w68, 
            w69=> c1_n21_w69, 
            w70=> c1_n21_w70, 
            w71=> c1_n21_w71, 
            w72=> c1_n21_w72, 
            w73=> c1_n21_w73, 
            w74=> c1_n21_w74, 
            w75=> c1_n21_w75, 
            w76=> c1_n21_w76, 
            w77=> c1_n21_w77, 
            w78=> c1_n21_w78, 
            w79=> c1_n21_w79, 
            w80=> c1_n21_w80, 
            w81=> c1_n21_w81, 
            w82=> c1_n21_w82, 
            w83=> c1_n21_w83, 
            w84=> c1_n21_w84, 
            w85=> c1_n21_w85, 
            w86=> c1_n21_w86, 
            w87=> c1_n21_w87, 
            w88=> c1_n21_w88, 
            w89=> c1_n21_w89, 
            w90=> c1_n21_w90, 
            w91=> c1_n21_w91, 
            w92=> c1_n21_w92, 
            w93=> c1_n21_w93, 
            w94=> c1_n21_w94, 
            w95=> c1_n21_w95, 
            w96=> c1_n21_w96, 
            w97=> c1_n21_w97, 
            w98=> c1_n21_w98, 
            w99=> c1_n21_w99, 
            w100=> c1_n21_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n21_y
   );           
            
neuron_inst_22: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n22_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n22_w1, 
            w2=> c1_n22_w2, 
            w3=> c1_n22_w3, 
            w4=> c1_n22_w4, 
            w5=> c1_n22_w5, 
            w6=> c1_n22_w6, 
            w7=> c1_n22_w7, 
            w8=> c1_n22_w8, 
            w9=> c1_n22_w9, 
            w10=> c1_n22_w10, 
            w11=> c1_n22_w11, 
            w12=> c1_n22_w12, 
            w13=> c1_n22_w13, 
            w14=> c1_n22_w14, 
            w15=> c1_n22_w15, 
            w16=> c1_n22_w16, 
            w17=> c1_n22_w17, 
            w18=> c1_n22_w18, 
            w19=> c1_n22_w19, 
            w20=> c1_n22_w20, 
            w21=> c1_n22_w21, 
            w22=> c1_n22_w22, 
            w23=> c1_n22_w23, 
            w24=> c1_n22_w24, 
            w25=> c1_n22_w25, 
            w26=> c1_n22_w26, 
            w27=> c1_n22_w27, 
            w28=> c1_n22_w28, 
            w29=> c1_n22_w29, 
            w30=> c1_n22_w30, 
            w31=> c1_n22_w31, 
            w32=> c1_n22_w32, 
            w33=> c1_n22_w33, 
            w34=> c1_n22_w34, 
            w35=> c1_n22_w35, 
            w36=> c1_n22_w36, 
            w37=> c1_n22_w37, 
            w38=> c1_n22_w38, 
            w39=> c1_n22_w39, 
            w40=> c1_n22_w40, 
            w41=> c1_n22_w41, 
            w42=> c1_n22_w42, 
            w43=> c1_n22_w43, 
            w44=> c1_n22_w44, 
            w45=> c1_n22_w45, 
            w46=> c1_n22_w46, 
            w47=> c1_n22_w47, 
            w48=> c1_n22_w48, 
            w49=> c1_n22_w49, 
            w50=> c1_n22_w50, 
            w51=> c1_n22_w51, 
            w52=> c1_n22_w52, 
            w53=> c1_n22_w53, 
            w54=> c1_n22_w54, 
            w55=> c1_n22_w55, 
            w56=> c1_n22_w56, 
            w57=> c1_n22_w57, 
            w58=> c1_n22_w58, 
            w59=> c1_n22_w59, 
            w60=> c1_n22_w60, 
            w61=> c1_n22_w61, 
            w62=> c1_n22_w62, 
            w63=> c1_n22_w63, 
            w64=> c1_n22_w64, 
            w65=> c1_n22_w65, 
            w66=> c1_n22_w66, 
            w67=> c1_n22_w67, 
            w68=> c1_n22_w68, 
            w69=> c1_n22_w69, 
            w70=> c1_n22_w70, 
            w71=> c1_n22_w71, 
            w72=> c1_n22_w72, 
            w73=> c1_n22_w73, 
            w74=> c1_n22_w74, 
            w75=> c1_n22_w75, 
            w76=> c1_n22_w76, 
            w77=> c1_n22_w77, 
            w78=> c1_n22_w78, 
            w79=> c1_n22_w79, 
            w80=> c1_n22_w80, 
            w81=> c1_n22_w81, 
            w82=> c1_n22_w82, 
            w83=> c1_n22_w83, 
            w84=> c1_n22_w84, 
            w85=> c1_n22_w85, 
            w86=> c1_n22_w86, 
            w87=> c1_n22_w87, 
            w88=> c1_n22_w88, 
            w89=> c1_n22_w89, 
            w90=> c1_n22_w90, 
            w91=> c1_n22_w91, 
            w92=> c1_n22_w92, 
            w93=> c1_n22_w93, 
            w94=> c1_n22_w94, 
            w95=> c1_n22_w95, 
            w96=> c1_n22_w96, 
            w97=> c1_n22_w97, 
            w98=> c1_n22_w98, 
            w99=> c1_n22_w99, 
            w100=> c1_n22_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n22_y
   );           
            
neuron_inst_23: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n23_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n23_w1, 
            w2=> c1_n23_w2, 
            w3=> c1_n23_w3, 
            w4=> c1_n23_w4, 
            w5=> c1_n23_w5, 
            w6=> c1_n23_w6, 
            w7=> c1_n23_w7, 
            w8=> c1_n23_w8, 
            w9=> c1_n23_w9, 
            w10=> c1_n23_w10, 
            w11=> c1_n23_w11, 
            w12=> c1_n23_w12, 
            w13=> c1_n23_w13, 
            w14=> c1_n23_w14, 
            w15=> c1_n23_w15, 
            w16=> c1_n23_w16, 
            w17=> c1_n23_w17, 
            w18=> c1_n23_w18, 
            w19=> c1_n23_w19, 
            w20=> c1_n23_w20, 
            w21=> c1_n23_w21, 
            w22=> c1_n23_w22, 
            w23=> c1_n23_w23, 
            w24=> c1_n23_w24, 
            w25=> c1_n23_w25, 
            w26=> c1_n23_w26, 
            w27=> c1_n23_w27, 
            w28=> c1_n23_w28, 
            w29=> c1_n23_w29, 
            w30=> c1_n23_w30, 
            w31=> c1_n23_w31, 
            w32=> c1_n23_w32, 
            w33=> c1_n23_w33, 
            w34=> c1_n23_w34, 
            w35=> c1_n23_w35, 
            w36=> c1_n23_w36, 
            w37=> c1_n23_w37, 
            w38=> c1_n23_w38, 
            w39=> c1_n23_w39, 
            w40=> c1_n23_w40, 
            w41=> c1_n23_w41, 
            w42=> c1_n23_w42, 
            w43=> c1_n23_w43, 
            w44=> c1_n23_w44, 
            w45=> c1_n23_w45, 
            w46=> c1_n23_w46, 
            w47=> c1_n23_w47, 
            w48=> c1_n23_w48, 
            w49=> c1_n23_w49, 
            w50=> c1_n23_w50, 
            w51=> c1_n23_w51, 
            w52=> c1_n23_w52, 
            w53=> c1_n23_w53, 
            w54=> c1_n23_w54, 
            w55=> c1_n23_w55, 
            w56=> c1_n23_w56, 
            w57=> c1_n23_w57, 
            w58=> c1_n23_w58, 
            w59=> c1_n23_w59, 
            w60=> c1_n23_w60, 
            w61=> c1_n23_w61, 
            w62=> c1_n23_w62, 
            w63=> c1_n23_w63, 
            w64=> c1_n23_w64, 
            w65=> c1_n23_w65, 
            w66=> c1_n23_w66, 
            w67=> c1_n23_w67, 
            w68=> c1_n23_w68, 
            w69=> c1_n23_w69, 
            w70=> c1_n23_w70, 
            w71=> c1_n23_w71, 
            w72=> c1_n23_w72, 
            w73=> c1_n23_w73, 
            w74=> c1_n23_w74, 
            w75=> c1_n23_w75, 
            w76=> c1_n23_w76, 
            w77=> c1_n23_w77, 
            w78=> c1_n23_w78, 
            w79=> c1_n23_w79, 
            w80=> c1_n23_w80, 
            w81=> c1_n23_w81, 
            w82=> c1_n23_w82, 
            w83=> c1_n23_w83, 
            w84=> c1_n23_w84, 
            w85=> c1_n23_w85, 
            w86=> c1_n23_w86, 
            w87=> c1_n23_w87, 
            w88=> c1_n23_w88, 
            w89=> c1_n23_w89, 
            w90=> c1_n23_w90, 
            w91=> c1_n23_w91, 
            w92=> c1_n23_w92, 
            w93=> c1_n23_w93, 
            w94=> c1_n23_w94, 
            w95=> c1_n23_w95, 
            w96=> c1_n23_w96, 
            w97=> c1_n23_w97, 
            w98=> c1_n23_w98, 
            w99=> c1_n23_w99, 
            w100=> c1_n23_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n23_y
   );           
            
neuron_inst_24: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n24_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n24_w1, 
            w2=> c1_n24_w2, 
            w3=> c1_n24_w3, 
            w4=> c1_n24_w4, 
            w5=> c1_n24_w5, 
            w6=> c1_n24_w6, 
            w7=> c1_n24_w7, 
            w8=> c1_n24_w8, 
            w9=> c1_n24_w9, 
            w10=> c1_n24_w10, 
            w11=> c1_n24_w11, 
            w12=> c1_n24_w12, 
            w13=> c1_n24_w13, 
            w14=> c1_n24_w14, 
            w15=> c1_n24_w15, 
            w16=> c1_n24_w16, 
            w17=> c1_n24_w17, 
            w18=> c1_n24_w18, 
            w19=> c1_n24_w19, 
            w20=> c1_n24_w20, 
            w21=> c1_n24_w21, 
            w22=> c1_n24_w22, 
            w23=> c1_n24_w23, 
            w24=> c1_n24_w24, 
            w25=> c1_n24_w25, 
            w26=> c1_n24_w26, 
            w27=> c1_n24_w27, 
            w28=> c1_n24_w28, 
            w29=> c1_n24_w29, 
            w30=> c1_n24_w30, 
            w31=> c1_n24_w31, 
            w32=> c1_n24_w32, 
            w33=> c1_n24_w33, 
            w34=> c1_n24_w34, 
            w35=> c1_n24_w35, 
            w36=> c1_n24_w36, 
            w37=> c1_n24_w37, 
            w38=> c1_n24_w38, 
            w39=> c1_n24_w39, 
            w40=> c1_n24_w40, 
            w41=> c1_n24_w41, 
            w42=> c1_n24_w42, 
            w43=> c1_n24_w43, 
            w44=> c1_n24_w44, 
            w45=> c1_n24_w45, 
            w46=> c1_n24_w46, 
            w47=> c1_n24_w47, 
            w48=> c1_n24_w48, 
            w49=> c1_n24_w49, 
            w50=> c1_n24_w50, 
            w51=> c1_n24_w51, 
            w52=> c1_n24_w52, 
            w53=> c1_n24_w53, 
            w54=> c1_n24_w54, 
            w55=> c1_n24_w55, 
            w56=> c1_n24_w56, 
            w57=> c1_n24_w57, 
            w58=> c1_n24_w58, 
            w59=> c1_n24_w59, 
            w60=> c1_n24_w60, 
            w61=> c1_n24_w61, 
            w62=> c1_n24_w62, 
            w63=> c1_n24_w63, 
            w64=> c1_n24_w64, 
            w65=> c1_n24_w65, 
            w66=> c1_n24_w66, 
            w67=> c1_n24_w67, 
            w68=> c1_n24_w68, 
            w69=> c1_n24_w69, 
            w70=> c1_n24_w70, 
            w71=> c1_n24_w71, 
            w72=> c1_n24_w72, 
            w73=> c1_n24_w73, 
            w74=> c1_n24_w74, 
            w75=> c1_n24_w75, 
            w76=> c1_n24_w76, 
            w77=> c1_n24_w77, 
            w78=> c1_n24_w78, 
            w79=> c1_n24_w79, 
            w80=> c1_n24_w80, 
            w81=> c1_n24_w81, 
            w82=> c1_n24_w82, 
            w83=> c1_n24_w83, 
            w84=> c1_n24_w84, 
            w85=> c1_n24_w85, 
            w86=> c1_n24_w86, 
            w87=> c1_n24_w87, 
            w88=> c1_n24_w88, 
            w89=> c1_n24_w89, 
            w90=> c1_n24_w90, 
            w91=> c1_n24_w91, 
            w92=> c1_n24_w92, 
            w93=> c1_n24_w93, 
            w94=> c1_n24_w94, 
            w95=> c1_n24_w95, 
            w96=> c1_n24_w96, 
            w97=> c1_n24_w97, 
            w98=> c1_n24_w98, 
            w99=> c1_n24_w99, 
            w100=> c1_n24_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n24_y
   );           
            
neuron_inst_25: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n25_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n25_w1, 
            w2=> c1_n25_w2, 
            w3=> c1_n25_w3, 
            w4=> c1_n25_w4, 
            w5=> c1_n25_w5, 
            w6=> c1_n25_w6, 
            w7=> c1_n25_w7, 
            w8=> c1_n25_w8, 
            w9=> c1_n25_w9, 
            w10=> c1_n25_w10, 
            w11=> c1_n25_w11, 
            w12=> c1_n25_w12, 
            w13=> c1_n25_w13, 
            w14=> c1_n25_w14, 
            w15=> c1_n25_w15, 
            w16=> c1_n25_w16, 
            w17=> c1_n25_w17, 
            w18=> c1_n25_w18, 
            w19=> c1_n25_w19, 
            w20=> c1_n25_w20, 
            w21=> c1_n25_w21, 
            w22=> c1_n25_w22, 
            w23=> c1_n25_w23, 
            w24=> c1_n25_w24, 
            w25=> c1_n25_w25, 
            w26=> c1_n25_w26, 
            w27=> c1_n25_w27, 
            w28=> c1_n25_w28, 
            w29=> c1_n25_w29, 
            w30=> c1_n25_w30, 
            w31=> c1_n25_w31, 
            w32=> c1_n25_w32, 
            w33=> c1_n25_w33, 
            w34=> c1_n25_w34, 
            w35=> c1_n25_w35, 
            w36=> c1_n25_w36, 
            w37=> c1_n25_w37, 
            w38=> c1_n25_w38, 
            w39=> c1_n25_w39, 
            w40=> c1_n25_w40, 
            w41=> c1_n25_w41, 
            w42=> c1_n25_w42, 
            w43=> c1_n25_w43, 
            w44=> c1_n25_w44, 
            w45=> c1_n25_w45, 
            w46=> c1_n25_w46, 
            w47=> c1_n25_w47, 
            w48=> c1_n25_w48, 
            w49=> c1_n25_w49, 
            w50=> c1_n25_w50, 
            w51=> c1_n25_w51, 
            w52=> c1_n25_w52, 
            w53=> c1_n25_w53, 
            w54=> c1_n25_w54, 
            w55=> c1_n25_w55, 
            w56=> c1_n25_w56, 
            w57=> c1_n25_w57, 
            w58=> c1_n25_w58, 
            w59=> c1_n25_w59, 
            w60=> c1_n25_w60, 
            w61=> c1_n25_w61, 
            w62=> c1_n25_w62, 
            w63=> c1_n25_w63, 
            w64=> c1_n25_w64, 
            w65=> c1_n25_w65, 
            w66=> c1_n25_w66, 
            w67=> c1_n25_w67, 
            w68=> c1_n25_w68, 
            w69=> c1_n25_w69, 
            w70=> c1_n25_w70, 
            w71=> c1_n25_w71, 
            w72=> c1_n25_w72, 
            w73=> c1_n25_w73, 
            w74=> c1_n25_w74, 
            w75=> c1_n25_w75, 
            w76=> c1_n25_w76, 
            w77=> c1_n25_w77, 
            w78=> c1_n25_w78, 
            w79=> c1_n25_w79, 
            w80=> c1_n25_w80, 
            w81=> c1_n25_w81, 
            w82=> c1_n25_w82, 
            w83=> c1_n25_w83, 
            w84=> c1_n25_w84, 
            w85=> c1_n25_w85, 
            w86=> c1_n25_w86, 
            w87=> c1_n25_w87, 
            w88=> c1_n25_w88, 
            w89=> c1_n25_w89, 
            w90=> c1_n25_w90, 
            w91=> c1_n25_w91, 
            w92=> c1_n25_w92, 
            w93=> c1_n25_w93, 
            w94=> c1_n25_w94, 
            w95=> c1_n25_w95, 
            w96=> c1_n25_w96, 
            w97=> c1_n25_w97, 
            w98=> c1_n25_w98, 
            w99=> c1_n25_w99, 
            w100=> c1_n25_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n25_y
   );           
            
neuron_inst_26: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n26_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n26_w1, 
            w2=> c1_n26_w2, 
            w3=> c1_n26_w3, 
            w4=> c1_n26_w4, 
            w5=> c1_n26_w5, 
            w6=> c1_n26_w6, 
            w7=> c1_n26_w7, 
            w8=> c1_n26_w8, 
            w9=> c1_n26_w9, 
            w10=> c1_n26_w10, 
            w11=> c1_n26_w11, 
            w12=> c1_n26_w12, 
            w13=> c1_n26_w13, 
            w14=> c1_n26_w14, 
            w15=> c1_n26_w15, 
            w16=> c1_n26_w16, 
            w17=> c1_n26_w17, 
            w18=> c1_n26_w18, 
            w19=> c1_n26_w19, 
            w20=> c1_n26_w20, 
            w21=> c1_n26_w21, 
            w22=> c1_n26_w22, 
            w23=> c1_n26_w23, 
            w24=> c1_n26_w24, 
            w25=> c1_n26_w25, 
            w26=> c1_n26_w26, 
            w27=> c1_n26_w27, 
            w28=> c1_n26_w28, 
            w29=> c1_n26_w29, 
            w30=> c1_n26_w30, 
            w31=> c1_n26_w31, 
            w32=> c1_n26_w32, 
            w33=> c1_n26_w33, 
            w34=> c1_n26_w34, 
            w35=> c1_n26_w35, 
            w36=> c1_n26_w36, 
            w37=> c1_n26_w37, 
            w38=> c1_n26_w38, 
            w39=> c1_n26_w39, 
            w40=> c1_n26_w40, 
            w41=> c1_n26_w41, 
            w42=> c1_n26_w42, 
            w43=> c1_n26_w43, 
            w44=> c1_n26_w44, 
            w45=> c1_n26_w45, 
            w46=> c1_n26_w46, 
            w47=> c1_n26_w47, 
            w48=> c1_n26_w48, 
            w49=> c1_n26_w49, 
            w50=> c1_n26_w50, 
            w51=> c1_n26_w51, 
            w52=> c1_n26_w52, 
            w53=> c1_n26_w53, 
            w54=> c1_n26_w54, 
            w55=> c1_n26_w55, 
            w56=> c1_n26_w56, 
            w57=> c1_n26_w57, 
            w58=> c1_n26_w58, 
            w59=> c1_n26_w59, 
            w60=> c1_n26_w60, 
            w61=> c1_n26_w61, 
            w62=> c1_n26_w62, 
            w63=> c1_n26_w63, 
            w64=> c1_n26_w64, 
            w65=> c1_n26_w65, 
            w66=> c1_n26_w66, 
            w67=> c1_n26_w67, 
            w68=> c1_n26_w68, 
            w69=> c1_n26_w69, 
            w70=> c1_n26_w70, 
            w71=> c1_n26_w71, 
            w72=> c1_n26_w72, 
            w73=> c1_n26_w73, 
            w74=> c1_n26_w74, 
            w75=> c1_n26_w75, 
            w76=> c1_n26_w76, 
            w77=> c1_n26_w77, 
            w78=> c1_n26_w78, 
            w79=> c1_n26_w79, 
            w80=> c1_n26_w80, 
            w81=> c1_n26_w81, 
            w82=> c1_n26_w82, 
            w83=> c1_n26_w83, 
            w84=> c1_n26_w84, 
            w85=> c1_n26_w85, 
            w86=> c1_n26_w86, 
            w87=> c1_n26_w87, 
            w88=> c1_n26_w88, 
            w89=> c1_n26_w89, 
            w90=> c1_n26_w90, 
            w91=> c1_n26_w91, 
            w92=> c1_n26_w92, 
            w93=> c1_n26_w93, 
            w94=> c1_n26_w94, 
            w95=> c1_n26_w95, 
            w96=> c1_n26_w96, 
            w97=> c1_n26_w97, 
            w98=> c1_n26_w98, 
            w99=> c1_n26_w99, 
            w100=> c1_n26_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n26_y
   );           
            
neuron_inst_27: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n27_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n27_w1, 
            w2=> c1_n27_w2, 
            w3=> c1_n27_w3, 
            w4=> c1_n27_w4, 
            w5=> c1_n27_w5, 
            w6=> c1_n27_w6, 
            w7=> c1_n27_w7, 
            w8=> c1_n27_w8, 
            w9=> c1_n27_w9, 
            w10=> c1_n27_w10, 
            w11=> c1_n27_w11, 
            w12=> c1_n27_w12, 
            w13=> c1_n27_w13, 
            w14=> c1_n27_w14, 
            w15=> c1_n27_w15, 
            w16=> c1_n27_w16, 
            w17=> c1_n27_w17, 
            w18=> c1_n27_w18, 
            w19=> c1_n27_w19, 
            w20=> c1_n27_w20, 
            w21=> c1_n27_w21, 
            w22=> c1_n27_w22, 
            w23=> c1_n27_w23, 
            w24=> c1_n27_w24, 
            w25=> c1_n27_w25, 
            w26=> c1_n27_w26, 
            w27=> c1_n27_w27, 
            w28=> c1_n27_w28, 
            w29=> c1_n27_w29, 
            w30=> c1_n27_w30, 
            w31=> c1_n27_w31, 
            w32=> c1_n27_w32, 
            w33=> c1_n27_w33, 
            w34=> c1_n27_w34, 
            w35=> c1_n27_w35, 
            w36=> c1_n27_w36, 
            w37=> c1_n27_w37, 
            w38=> c1_n27_w38, 
            w39=> c1_n27_w39, 
            w40=> c1_n27_w40, 
            w41=> c1_n27_w41, 
            w42=> c1_n27_w42, 
            w43=> c1_n27_w43, 
            w44=> c1_n27_w44, 
            w45=> c1_n27_w45, 
            w46=> c1_n27_w46, 
            w47=> c1_n27_w47, 
            w48=> c1_n27_w48, 
            w49=> c1_n27_w49, 
            w50=> c1_n27_w50, 
            w51=> c1_n27_w51, 
            w52=> c1_n27_w52, 
            w53=> c1_n27_w53, 
            w54=> c1_n27_w54, 
            w55=> c1_n27_w55, 
            w56=> c1_n27_w56, 
            w57=> c1_n27_w57, 
            w58=> c1_n27_w58, 
            w59=> c1_n27_w59, 
            w60=> c1_n27_w60, 
            w61=> c1_n27_w61, 
            w62=> c1_n27_w62, 
            w63=> c1_n27_w63, 
            w64=> c1_n27_w64, 
            w65=> c1_n27_w65, 
            w66=> c1_n27_w66, 
            w67=> c1_n27_w67, 
            w68=> c1_n27_w68, 
            w69=> c1_n27_w69, 
            w70=> c1_n27_w70, 
            w71=> c1_n27_w71, 
            w72=> c1_n27_w72, 
            w73=> c1_n27_w73, 
            w74=> c1_n27_w74, 
            w75=> c1_n27_w75, 
            w76=> c1_n27_w76, 
            w77=> c1_n27_w77, 
            w78=> c1_n27_w78, 
            w79=> c1_n27_w79, 
            w80=> c1_n27_w80, 
            w81=> c1_n27_w81, 
            w82=> c1_n27_w82, 
            w83=> c1_n27_w83, 
            w84=> c1_n27_w84, 
            w85=> c1_n27_w85, 
            w86=> c1_n27_w86, 
            w87=> c1_n27_w87, 
            w88=> c1_n27_w88, 
            w89=> c1_n27_w89, 
            w90=> c1_n27_w90, 
            w91=> c1_n27_w91, 
            w92=> c1_n27_w92, 
            w93=> c1_n27_w93, 
            w94=> c1_n27_w94, 
            w95=> c1_n27_w95, 
            w96=> c1_n27_w96, 
            w97=> c1_n27_w97, 
            w98=> c1_n27_w98, 
            w99=> c1_n27_w99, 
            w100=> c1_n27_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n27_y
   );           
            
neuron_inst_28: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n28_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n28_w1, 
            w2=> c1_n28_w2, 
            w3=> c1_n28_w3, 
            w4=> c1_n28_w4, 
            w5=> c1_n28_w5, 
            w6=> c1_n28_w6, 
            w7=> c1_n28_w7, 
            w8=> c1_n28_w8, 
            w9=> c1_n28_w9, 
            w10=> c1_n28_w10, 
            w11=> c1_n28_w11, 
            w12=> c1_n28_w12, 
            w13=> c1_n28_w13, 
            w14=> c1_n28_w14, 
            w15=> c1_n28_w15, 
            w16=> c1_n28_w16, 
            w17=> c1_n28_w17, 
            w18=> c1_n28_w18, 
            w19=> c1_n28_w19, 
            w20=> c1_n28_w20, 
            w21=> c1_n28_w21, 
            w22=> c1_n28_w22, 
            w23=> c1_n28_w23, 
            w24=> c1_n28_w24, 
            w25=> c1_n28_w25, 
            w26=> c1_n28_w26, 
            w27=> c1_n28_w27, 
            w28=> c1_n28_w28, 
            w29=> c1_n28_w29, 
            w30=> c1_n28_w30, 
            w31=> c1_n28_w31, 
            w32=> c1_n28_w32, 
            w33=> c1_n28_w33, 
            w34=> c1_n28_w34, 
            w35=> c1_n28_w35, 
            w36=> c1_n28_w36, 
            w37=> c1_n28_w37, 
            w38=> c1_n28_w38, 
            w39=> c1_n28_w39, 
            w40=> c1_n28_w40, 
            w41=> c1_n28_w41, 
            w42=> c1_n28_w42, 
            w43=> c1_n28_w43, 
            w44=> c1_n28_w44, 
            w45=> c1_n28_w45, 
            w46=> c1_n28_w46, 
            w47=> c1_n28_w47, 
            w48=> c1_n28_w48, 
            w49=> c1_n28_w49, 
            w50=> c1_n28_w50, 
            w51=> c1_n28_w51, 
            w52=> c1_n28_w52, 
            w53=> c1_n28_w53, 
            w54=> c1_n28_w54, 
            w55=> c1_n28_w55, 
            w56=> c1_n28_w56, 
            w57=> c1_n28_w57, 
            w58=> c1_n28_w58, 
            w59=> c1_n28_w59, 
            w60=> c1_n28_w60, 
            w61=> c1_n28_w61, 
            w62=> c1_n28_w62, 
            w63=> c1_n28_w63, 
            w64=> c1_n28_w64, 
            w65=> c1_n28_w65, 
            w66=> c1_n28_w66, 
            w67=> c1_n28_w67, 
            w68=> c1_n28_w68, 
            w69=> c1_n28_w69, 
            w70=> c1_n28_w70, 
            w71=> c1_n28_w71, 
            w72=> c1_n28_w72, 
            w73=> c1_n28_w73, 
            w74=> c1_n28_w74, 
            w75=> c1_n28_w75, 
            w76=> c1_n28_w76, 
            w77=> c1_n28_w77, 
            w78=> c1_n28_w78, 
            w79=> c1_n28_w79, 
            w80=> c1_n28_w80, 
            w81=> c1_n28_w81, 
            w82=> c1_n28_w82, 
            w83=> c1_n28_w83, 
            w84=> c1_n28_w84, 
            w85=> c1_n28_w85, 
            w86=> c1_n28_w86, 
            w87=> c1_n28_w87, 
            w88=> c1_n28_w88, 
            w89=> c1_n28_w89, 
            w90=> c1_n28_w90, 
            w91=> c1_n28_w91, 
            w92=> c1_n28_w92, 
            w93=> c1_n28_w93, 
            w94=> c1_n28_w94, 
            w95=> c1_n28_w95, 
            w96=> c1_n28_w96, 
            w97=> c1_n28_w97, 
            w98=> c1_n28_w98, 
            w99=> c1_n28_w99, 
            w100=> c1_n28_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n28_y
   );           
            
neuron_inst_29: ENTITY work.neuron_comb_Barriers_Leaky_ReLU_100n_8bit_mul0_add0_v0_v0_unsigned
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            -- ['IN']['SIGNED'] 
            bias=> c1_n29_bias, 
            -- ['IN']['SIGNED_num_inputs'] 
            x1=> x1, 
            x2=> x2, 
            x3=> x3, 
            x4=> x4, 
            x5=> x5, 
            x6=> x6, 
            x7=> x7, 
            x8=> x8, 
            x9=> x9, 
            x10=> x10, 
            x11=> x11, 
            x12=> x12, 
            x13=> x13, 
            x14=> x14, 
            x15=> x15, 
            x16=> x16, 
            x17=> x17, 
            x18=> x18, 
            x19=> x19, 
            x20=> x20, 
            x21=> x21, 
            x22=> x22, 
            x23=> x23, 
            x24=> x24, 
            x25=> x25, 
            x26=> x26, 
            x27=> x27, 
            x28=> x28, 
            x29=> x29, 
            x30=> x30, 
            x31=> x31, 
            x32=> x32, 
            x33=> x33, 
            x34=> x34, 
            x35=> x35, 
            x36=> x36, 
            x37=> x37, 
            x38=> x38, 
            x39=> x39, 
            x40=> x40, 
            x41=> x41, 
            x42=> x42, 
            x43=> x43, 
            x44=> x44, 
            x45=> x45, 
            x46=> x46, 
            x47=> x47, 
            x48=> x48, 
            x49=> x49, 
            x50=> x50, 
            x51=> x51, 
            x52=> x52, 
            x53=> x53, 
            x54=> x54, 
            x55=> x55, 
            x56=> x56, 
            x57=> x57, 
            x58=> x58, 
            x59=> x59, 
            x60=> x60, 
            x61=> x61, 
            x62=> x62, 
            x63=> x63, 
            x64=> x64, 
            x65=> x65, 
            x66=> x66, 
            x67=> x67, 
            x68=> x68, 
            x69=> x69, 
            x70=> x70, 
            x71=> x71, 
            x72=> x72, 
            x73=> x73, 
            x74=> x74, 
            x75=> x75, 
            x76=> x76, 
            x77=> x77, 
            x78=> x78, 
            x79=> x79, 
            x80=> x80, 
            x81=> x81, 
            x82=> x82, 
            x83=> x83, 
            x84=> x84, 
            x85=> x85, 
            x86=> x86, 
            x87=> x87, 
            x88=> x88, 
            x89=> x89, 
            x90=> x90, 
            x91=> x91, 
            x92=> x92, 
            x93=> x93, 
            x94=> x94, 
            x95=> x95, 
            x96=> x96, 
            x97=> x97, 
            x98=> x98, 
            x99=> x99, 
            x100=> x100, 
            w1=> c1_n29_w1, 
            w2=> c1_n29_w2, 
            w3=> c1_n29_w3, 
            w4=> c1_n29_w4, 
            w5=> c1_n29_w5, 
            w6=> c1_n29_w6, 
            w7=> c1_n29_w7, 
            w8=> c1_n29_w8, 
            w9=> c1_n29_w9, 
            w10=> c1_n29_w10, 
            w11=> c1_n29_w11, 
            w12=> c1_n29_w12, 
            w13=> c1_n29_w13, 
            w14=> c1_n29_w14, 
            w15=> c1_n29_w15, 
            w16=> c1_n29_w16, 
            w17=> c1_n29_w17, 
            w18=> c1_n29_w18, 
            w19=> c1_n29_w19, 
            w20=> c1_n29_w20, 
            w21=> c1_n29_w21, 
            w22=> c1_n29_w22, 
            w23=> c1_n29_w23, 
            w24=> c1_n29_w24, 
            w25=> c1_n29_w25, 
            w26=> c1_n29_w26, 
            w27=> c1_n29_w27, 
            w28=> c1_n29_w28, 
            w29=> c1_n29_w29, 
            w30=> c1_n29_w30, 
            w31=> c1_n29_w31, 
            w32=> c1_n29_w32, 
            w33=> c1_n29_w33, 
            w34=> c1_n29_w34, 
            w35=> c1_n29_w35, 
            w36=> c1_n29_w36, 
            w37=> c1_n29_w37, 
            w38=> c1_n29_w38, 
            w39=> c1_n29_w39, 
            w40=> c1_n29_w40, 
            w41=> c1_n29_w41, 
            w42=> c1_n29_w42, 
            w43=> c1_n29_w43, 
            w44=> c1_n29_w44, 
            w45=> c1_n29_w45, 
            w46=> c1_n29_w46, 
            w47=> c1_n29_w47, 
            w48=> c1_n29_w48, 
            w49=> c1_n29_w49, 
            w50=> c1_n29_w50, 
            w51=> c1_n29_w51, 
            w52=> c1_n29_w52, 
            w53=> c1_n29_w53, 
            w54=> c1_n29_w54, 
            w55=> c1_n29_w55, 
            w56=> c1_n29_w56, 
            w57=> c1_n29_w57, 
            w58=> c1_n29_w58, 
            w59=> c1_n29_w59, 
            w60=> c1_n29_w60, 
            w61=> c1_n29_w61, 
            w62=> c1_n29_w62, 
            w63=> c1_n29_w63, 
            w64=> c1_n29_w64, 
            w65=> c1_n29_w65, 
            w66=> c1_n29_w66, 
            w67=> c1_n29_w67, 
            w68=> c1_n29_w68, 
            w69=> c1_n29_w69, 
            w70=> c1_n29_w70, 
            w71=> c1_n29_w71, 
            w72=> c1_n29_w72, 
            w73=> c1_n29_w73, 
            w74=> c1_n29_w74, 
            w75=> c1_n29_w75, 
            w76=> c1_n29_w76, 
            w77=> c1_n29_w77, 
            w78=> c1_n29_w78, 
            w79=> c1_n29_w79, 
            w80=> c1_n29_w80, 
            w81=> c1_n29_w81, 
            w82=> c1_n29_w82, 
            w83=> c1_n29_w83, 
            w84=> c1_n29_w84, 
            w85=> c1_n29_w85, 
            w86=> c1_n29_w86, 
            w87=> c1_n29_w87, 
            w88=> c1_n29_w88, 
            w89=> c1_n29_w89, 
            w90=> c1_n29_w90, 
            w91=> c1_n29_w91, 
            w92=> c1_n29_w92, 
            w93=> c1_n29_w93, 
            w94=> c1_n29_w94, 
            w95=> c1_n29_w95, 
            w96=> c1_n29_w96, 
            w97=> c1_n29_w97, 
            w98=> c1_n29_w98, 
            w99=> c1_n29_w99, 
            w100=> c1_n29_w100, 
            ---------- Saidas ---------- 
            -- ['OUT']['SIGNED'] 
            y=> c1_n29_y
   );           
             
END ARCHITECTURE;
