LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.parameters.ALL;

ENTITY autoencoder_camada0_ReLU_5neuron_8bits_5n_signed IS
   GENERIC (
      BITS       : NATURAL := BITS;
      NUM_INPUTS : NATURAL := 5;
      TOTAL_BITS : NATURAL := 40
   );
   PORT (
      clk, rst, update_weights                                             : IN STD_LOGIC;
      -- IO_in: IN signed(TOTAL_BITS - 1 DOWNTO 0);
      IO_in                                                                : IN signed(TOTAL_BITS * NUM_INPUTS - 1 DOWNTO 0); -- todo
      c0_n0_W_in, c0_n1_W_in, c0_n2_W_in, c0_n3_W_in, c0_n4_W_in           : IN signed(BITS - 1 DOWNTO 0);
      ----------------------------------------------
      c0_n0_IO_out, c0_n1_IO_out, c0_n2_IO_out, c0_n3_IO_out, c0_n4_IO_out : OUT signed(BITS - 1 DOWNTO 0);
      c0_n0_W_out, c0_n1_W_out, c0_n2_W_out, c0_n3_W_out                   : OUT signed(BITS - 1 DOWNTO 0)
   );
END ENTITY;

ARCHITECTURE arch OF autoencoder_camada0_ReLU_5neuron_8bits_5n_signed IS
BEGIN

   neuron_inst_0 : ENTITY work.neuron_comb_ReLU_5n_8bit_signed_mult0_v0_add0_v0_out
      PORT MAP(
         ---------- Entradas ----------
         -- ['IN']['STD_LOGIC'] 
         clk            => clk,
         rst            => rst,
         update_weights => update_weights,
         -- ['IN']['manual'] 
         IO_in          => IO_in((TOTAL_BITS * 1) - 1 DOWNTO (TOTAL_BITS * 0)), -- todo
         W_in           => c0_n0_W_in,
         ---------- Saidas ----------
         -- ['OUT']['SIGNED'] 
         IO_out         => c0_n0_IO_out,
         -- ['OUT']['manual'] 
         W_out          => c0_n0_W_out
      );

   neuron_inst_1 : ENTITY work.neuron_comb_ReLU_5n_8bit_signed_mult0_v0_add0_v0_out
      PORT MAP(
         ---------- Entradas ----------
         -- ['IN']['STD_LOGIC'] 
         clk            => clk,
         rst            => rst,
         update_weights => update_weights,
         -- ['IN']['manual'] 
         IO_in          => IO_in((TOTAL_BITS * 2) - 1 DOWNTO (TOTAL_BITS * 1)), -- todo
         W_in           => c0_n1_W_in,
         ---------- Saidas ----------
         -- ['OUT']['SIGNED'] 
         IO_out         => c0_n1_IO_out,
         -- ['OUT']['manual'] 
         W_out          => c0_n1_W_out
      );

   neuron_inst_2 : ENTITY work.neuron_comb_ReLU_5n_8bit_signed_mult0_v0_add0_v0_out
      PORT MAP(
         ---------- Entradas ----------
         -- ['IN']['STD_LOGIC'] 
         clk            => clk,
         rst            => rst,
         update_weights => update_weights,
         -- ['IN']['manual'] 
         IO_in          => IO_in((TOTAL_BITS * 3) - 1 DOWNTO (TOTAL_BITS * 2)), -- todo
         W_in           => c0_n2_W_in,
         ---------- Saidas ----------
         -- ['OUT']['SIGNED'] 
         IO_out         => c0_n2_IO_out,
         -- ['OUT']['manual'] 
         W_out          => c0_n2_W_out
      );

   neuron_inst_3 : ENTITY work.neuron_comb_ReLU_5n_8bit_signed_mult0_v0_add0_v0_out
      PORT MAP(
         ---------- Entradas ----------
         -- ['IN']['STD_LOGIC'] 
         clk            => clk,
         rst            => rst,
         update_weights => update_weights,
         -- ['IN']['manual'] 
         IO_in          => IO_in((TOTAL_BITS * 4) - 1 DOWNTO (TOTAL_BITS * 3)), -- todo
         W_in           => c0_n3_W_in,
         ---------- Saidas ----------
         -- ['OUT']['SIGNED'] 
         IO_out         => c0_n3_IO_out,
         -- ['OUT']['manual'] 
         W_out          => c0_n3_W_out
      );

   neuron_inst_4 : ENTITY work.neuron_comb_ReLU_5n_8bit_signed_mult0_v0_add0_v0
      PORT MAP(
         ---------- Entradas ----------
         -- ['IN']['STD_LOGIC'] 
         clk            => clk,
         rst            => rst,
         update_weights => update_weights,
         -- ['IN']['manual'] 
         IO_in          => IO_in((TOTAL_BITS * 5) - 1 DOWNTO (TOTAL_BITS * 4)), -- todo
         W_in           => c0_n4_W_in,
         ---------- Saidas ----------
         -- ['OUT']['SIGNED'] 
         IO_out         => c0_n4_IO_out
      );

END ARCHITECTURE;