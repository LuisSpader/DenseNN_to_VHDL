LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.parameters.ALL;

  ENTITY  top IS
  GENERIC (
    BITS : NATURAL := BITS;
    NUM_INPUTS : NATURAL := 784;
    TOTAL_BITS : NATURAL := 6272
  );
  PORT (
      clk, rst, update_weights: IN STD_LOGIC;
      IO_in: IN signed(TOTAL_BITS - 1 DOWNTO 0);
      c0_n0_W_in, c0_n1_W_in, c0_n2_W_in, c0_n3_W_in, c0_n4_W_in, c0_n5_W_in, c0_n6_W_in, c0_n7_W_in, c0_n8_W_in, c0_n9_W_in, c0_n10_W_in, c0_n11_W_in, c0_n12_W_in, c0_n13_W_in, c0_n14_W_in, c0_n15_W_in, c0_n16_W_in, c0_n17_W_in, c0_n18_W_in, c0_n19_W_in, c0_n20_W_in, c0_n21_W_in, c0_n22_W_in, c0_n23_W_in, c0_n24_W_in, c0_n25_W_in, c0_n26_W_in, c0_n27_W_in, c0_n28_W_in, c0_n29_W_in, c0_n30_W_in, c0_n31_W_in, c0_n32_W_in, c0_n33_W_in, c0_n34_W_in, c0_n35_W_in, c0_n36_W_in, c0_n37_W_in, c0_n38_W_in, c0_n39_W_in, c0_n40_W_in, c0_n41_W_in, c0_n42_W_in, c0_n43_W_in, c0_n44_W_in, c0_n45_W_in, c0_n46_W_in, c0_n47_W_in, c0_n48_W_in, c0_n49_W_in, c0_n50_W_in, c0_n51_W_in, c0_n52_W_in, c0_n53_W_in, c0_n54_W_in, c0_n55_W_in, c0_n56_W_in, c0_n57_W_in, c0_n58_W_in, c0_n59_W_in, c0_n60_W_in, c0_n61_W_in, c0_n62_W_in, c0_n63_W_in, c0_n64_W_in, c0_n65_W_in, c0_n66_W_in, c0_n67_W_in, c0_n68_W_in, c0_n69_W_in, c0_n70_W_in, c0_n71_W_in, c0_n72_W_in, c0_n73_W_in, c0_n74_W_in, c0_n75_W_in, c0_n76_W_in, c0_n77_W_in, c0_n78_W_in, c0_n79_W_in, c0_n80_W_in, c0_n81_W_in, c0_n82_W_in, c0_n83_W_in, c0_n84_W_in, c0_n85_W_in, c0_n86_W_in, c0_n87_W_in, c0_n88_W_in, c0_n89_W_in, c0_n90_W_in, c0_n91_W_in, c0_n92_W_in, c0_n93_W_in, c0_n94_W_in, c0_n95_W_in, c0_n96_W_in, c0_n97_W_in, c0_n98_W_in, c0_n99_W_in, c0_n100_W_in, c0_n101_W_in, c0_n102_W_in, c0_n103_W_in, c0_n104_W_in, c0_n105_W_in, c0_n106_W_in, c0_n107_W_in, c0_n108_W_in, c0_n109_W_in, c0_n110_W_in, c0_n111_W_in, c0_n112_W_in, c0_n113_W_in, c0_n114_W_in, c0_n115_W_in, c0_n116_W_in, c0_n117_W_in, c0_n118_W_in, c0_n119_W_in, c0_n120_W_in, c0_n121_W_in, c0_n122_W_in, c0_n123_W_in, c0_n124_W_in, c0_n125_W_in, c0_n126_W_in, c0_n127_W_in: IN signed(BITS - 1 DOWNTO 0);
      ----------------------------------------------
      c6_n0_IO_out, c6_n1_IO_out, c6_n2_IO_out, c6_n3_IO_out, c6_n4_IO_out, c6_n5_IO_out, c6_n6_IO_out, c6_n7_IO_out, c6_n8_IO_out, c6_n9_IO_out, c6_n10_IO_out, c6_n11_IO_out, c6_n12_IO_out, c6_n13_IO_out, c6_n14_IO_out, c6_n15_IO_out, c6_n16_IO_out, c6_n17_IO_out, c6_n18_IO_out, c6_n19_IO_out, c6_n20_IO_out, c6_n21_IO_out, c6_n22_IO_out, c6_n23_IO_out, c6_n24_IO_out, c6_n25_IO_out, c6_n26_IO_out, c6_n27_IO_out, c6_n28_IO_out, c6_n29_IO_out, c6_n30_IO_out, c6_n31_IO_out, c6_n32_IO_out, c6_n33_IO_out, c6_n34_IO_out, c6_n35_IO_out, c6_n36_IO_out, c6_n37_IO_out, c6_n38_IO_out, c6_n39_IO_out, c6_n40_IO_out, c6_n41_IO_out, c6_n42_IO_out, c6_n43_IO_out, c6_n44_IO_out, c6_n45_IO_out, c6_n46_IO_out, c6_n47_IO_out, c6_n48_IO_out, c6_n49_IO_out, c6_n50_IO_out, c6_n51_IO_out, c6_n52_IO_out, c6_n53_IO_out, c6_n54_IO_out, c6_n55_IO_out, c6_n56_IO_out, c6_n57_IO_out, c6_n58_IO_out, c6_n59_IO_out, c6_n60_IO_out, c6_n61_IO_out, c6_n62_IO_out, c6_n63_IO_out, c6_n64_IO_out, c6_n65_IO_out, c6_n66_IO_out, c6_n67_IO_out, c6_n68_IO_out, c6_n69_IO_out, c6_n70_IO_out, c6_n71_IO_out, c6_n72_IO_out, c6_n73_IO_out, c6_n74_IO_out, c6_n75_IO_out, c6_n76_IO_out, c6_n77_IO_out, c6_n78_IO_out, c6_n79_IO_out, c6_n80_IO_out, c6_n81_IO_out, c6_n82_IO_out, c6_n83_IO_out, c6_n84_IO_out, c6_n85_IO_out, c6_n86_IO_out, c6_n87_IO_out, c6_n88_IO_out, c6_n89_IO_out, c6_n90_IO_out, c6_n91_IO_out, c6_n92_IO_out, c6_n93_IO_out, c6_n94_IO_out, c6_n95_IO_out, c6_n96_IO_out, c6_n97_IO_out, c6_n98_IO_out, c6_n99_IO_out, c6_n100_IO_out, c6_n101_IO_out, c6_n102_IO_out, c6_n103_IO_out, c6_n104_IO_out, c6_n105_IO_out, c6_n106_IO_out, c6_n107_IO_out, c6_n108_IO_out, c6_n109_IO_out, c6_n110_IO_out, c6_n111_IO_out, c6_n112_IO_out, c6_n113_IO_out, c6_n114_IO_out, c6_n115_IO_out, c6_n116_IO_out, c6_n117_IO_out, c6_n118_IO_out, c6_n119_IO_out, c6_n120_IO_out, c6_n121_IO_out, c6_n122_IO_out, c6_n123_IO_out, c6_n124_IO_out, c6_n125_IO_out, c6_n126_IO_out, c6_n127_IO_out: OUT signed(7 DOWNTO 0)
  );
  end ENTITY;

ARCHITECTURE arch OF  top  IS
-- SIGNALS
  SIGNAL c0_n0_W_out, c0_n1_W_out, c0_n2_W_out, c0_n3_W_out, c0_n4_W_out, c0_n5_W_out, c0_n6_W_out, c0_n7_W_out, c0_n8_W_out, c0_n9_W_out, c0_n10_W_out, c0_n11_W_out, c0_n12_W_out, c0_n13_W_out, c0_n14_W_out, c0_n15_W_out, c0_n16_W_out, c0_n17_W_out, c0_n18_W_out, c0_n19_W_out, c0_n20_W_out, c0_n21_W_out, c0_n22_W_out, c0_n23_W_out, c0_n24_W_out, c0_n25_W_out, c0_n26_W_out, c0_n27_W_out, c0_n28_W_out, c0_n29_W_out, c0_n30_W_out, c0_n31_W_out, c0_n32_W_out, c0_n33_W_out, c0_n34_W_out, c0_n35_W_out, c0_n36_W_out, c0_n37_W_out, c0_n38_W_out, c0_n39_W_out, c0_n40_W_out, c0_n41_W_out, c0_n42_W_out, c0_n43_W_out, c0_n44_W_out, c0_n45_W_out, c0_n46_W_out, c0_n47_W_out, c0_n48_W_out, c0_n49_W_out, c0_n50_W_out, c0_n51_W_out, c0_n52_W_out, c0_n53_W_out, c0_n54_W_out, c0_n55_W_out, c0_n56_W_out, c0_n57_W_out, c0_n58_W_out, c0_n59_W_out, c0_n60_W_out, c0_n61_W_out, c0_n62_W_out, c0_n63_W_out, c0_n64_W_out, c0_n65_W_out, c0_n66_W_out, c0_n67_W_out, c0_n68_W_out, c0_n69_W_out, c0_n70_W_out, c0_n71_W_out, c0_n72_W_out, c0_n73_W_out, c0_n74_W_out, c0_n75_W_out, c0_n76_W_out, c0_n77_W_out, c0_n78_W_out, c0_n79_W_out, c0_n80_W_out, c0_n81_W_out, c0_n82_W_out, c0_n83_W_out, c0_n84_W_out, c0_n85_W_out, c0_n86_W_out, c0_n87_W_out, c0_n88_W_out, c0_n89_W_out, c0_n90_W_out, c0_n91_W_out, c0_n92_W_out, c0_n93_W_out, c0_n94_W_out, c0_n95_W_out, c0_n96_W_out, c0_n97_W_out, c0_n98_W_out, c0_n99_W_out, c0_n100_W_out, c0_n101_W_out, c0_n102_W_out, c0_n103_W_out, c0_n104_W_out, c0_n105_W_out, c0_n106_W_out, c0_n107_W_out, c0_n108_W_out, c0_n109_W_out, c0_n110_W_out, c0_n111_W_out, c0_n112_W_out, c0_n113_W_out, c0_n114_W_out, c0_n115_W_out, c0_n116_W_out, c0_n117_W_out, c0_n118_W_out, c0_n119_W_out, c0_n120_W_out, c0_n121_W_out, c0_n122_W_out, c0_n123_W_out, c0_n124_W_out, c0_n125_W_out, c0_n126_W_out, c0_n127_W_out, c1_n0_W_out, c1_n1_W_out, c1_n2_W_out, c1_n3_W_out, c1_n4_W_out, c1_n5_W_out, c1_n6_W_out, c1_n7_W_out, c1_n8_W_out, c1_n9_W_out, c1_n10_W_out, c1_n11_W_out, c1_n12_W_out, c1_n13_W_out, c1_n14_W_out, c1_n15_W_out, c1_n16_W_out, c1_n17_W_out, c1_n18_W_out, c1_n19_W_out, c1_n20_W_out, c1_n21_W_out, c1_n22_W_out, c1_n23_W_out, c1_n24_W_out, c1_n25_W_out, c1_n26_W_out, c1_n27_W_out, c1_n28_W_out, c1_n29_W_out, c1_n30_W_out, c1_n31_W_out, c1_n32_W_out, c1_n33_W_out, c1_n34_W_out, c1_n35_W_out, c1_n36_W_out, c1_n37_W_out, c1_n38_W_out, c1_n39_W_out, c1_n40_W_out, c1_n41_W_out, c1_n42_W_out, c1_n43_W_out, c1_n44_W_out, c1_n45_W_out, c1_n46_W_out, c1_n47_W_out, c1_n48_W_out, c1_n49_W_out, c1_n50_W_out, c1_n51_W_out, c1_n52_W_out, c1_n53_W_out, c1_n54_W_out, c1_n55_W_out, c1_n56_W_out, c1_n57_W_out, c1_n58_W_out, c1_n59_W_out, c1_n60_W_out, c1_n61_W_out, c1_n62_W_out, c1_n63_W_out, c2_n0_W_out, c2_n1_W_out, c2_n2_W_out, c2_n3_W_out, c2_n4_W_out, c2_n5_W_out, c2_n6_W_out, c2_n7_W_out, c2_n8_W_out, c2_n9_W_out, c2_n10_W_out, c2_n11_W_out, c2_n12_W_out, c2_n13_W_out, c2_n14_W_out, c2_n15_W_out, c2_n16_W_out, c2_n17_W_out, c2_n18_W_out, c2_n19_W_out, c2_n20_W_out, c2_n21_W_out, c2_n22_W_out, c2_n23_W_out, c2_n24_W_out, c2_n25_W_out, c2_n26_W_out, c2_n27_W_out, c2_n28_W_out, c2_n29_W_out, c2_n30_W_out, c2_n31_W_out, c5_n32_W_out, c5_n33_W_out, c5_n34_W_out, c5_n35_W_out, c5_n36_W_out, c5_n37_W_out, c5_n38_W_out, c5_n39_W_out, c5_n40_W_out, c5_n41_W_out, c5_n42_W_out, c5_n43_W_out, c5_n44_W_out, c5_n45_W_out, c5_n46_W_out, c5_n47_W_out, c5_n48_W_out, c5_n49_W_out, c5_n50_W_out, c5_n51_W_out, c5_n52_W_out, c5_n53_W_out, c5_n54_W_out, c5_n55_W_out, c5_n56_W_out, c5_n57_W_out, c5_n58_W_out, c5_n59_W_out, c5_n60_W_out, c5_n61_W_out, c5_n62_W_out, c5_n63_W_out, c3_n0_W_out, c3_n1_W_out, c3_n2_W_out, c3_n3_W_out, c3_n4_W_out, c3_n5_W_out, c3_n6_W_out, c3_n7_W_out, c3_n8_W_out, c3_n9_W_out, c3_n10_W_out, c3_n11_W_out, c3_n12_W_out, c3_n13_W_out, c3_n14_W_out, c3_n15_W_out, c4_n16_W_out, c4_n17_W_out, c4_n18_W_out, c4_n19_W_out, c4_n20_W_out, c4_n21_W_out, c4_n22_W_out, c4_n23_W_out, c4_n24_W_out, c4_n25_W_out, c4_n26_W_out, c4_n27_W_out, c4_n28_W_out, c4_n29_W_out, c4_n30_W_out, c4_n31_W_out, c4_n0_W_out, c4_n1_W_out, c4_n2_W_out, c4_n3_W_out, c4_n4_W_out, c4_n5_W_out, c4_n6_W_out, c4_n7_W_out, c4_n8_W_out, c4_n9_W_out, c4_n10_W_out, c4_n11_W_out, c4_n12_W_out, c4_n13_W_out, c4_n14_W_out, c4_n15_W_out, c5_n16_W_out, c5_n17_W_out, c5_n18_W_out, c5_n19_W_out, c5_n20_W_out, c5_n21_W_out, c5_n22_W_out, c5_n23_W_out, c5_n24_W_out, c5_n25_W_out, c5_n26_W_out, c5_n27_W_out, c5_n28_W_out, c5_n29_W_out, c5_n30_W_out, c5_n31_W_out, c5_n0_W_out, c5_n1_W_out, c5_n2_W_out, c5_n3_W_out, c5_n4_W_out, c5_n5_W_out, c5_n6_W_out, c5_n7_W_out, c5_n8_W_out, c5_n9_W_out, c5_n10_W_out, c5_n11_W_out, c5_n12_W_out, c5_n13_W_out, c5_n14_W_out, c5_n15_W_out: signed(BITS - 1 DOWNTO 0);
  SIGNAL c1_IO_in:  signed((BITS*128) - 1 DOWNTO 0);
  SIGNAL c2_IO_in:  signed((BITS*64) - 1 DOWNTO 0);
  SIGNAL c3_IO_in:  signed((BITS*32) - 1 DOWNTO 0);
  SIGNAL c4_IO_in:  signed((BITS*16) - 1 DOWNTO 0);
  SIGNAL c5_IO_in:  signed((BITS*32) - 1 DOWNTO 0);
  SIGNAL c6_IO_in:  signed((BITS*64) - 1 DOWNTO 0);
  SIGNAL c0_n0_IO_out, c0_n1_IO_out, c0_n2_IO_out, c0_n3_IO_out, c0_n4_IO_out, c0_n5_IO_out, c0_n6_IO_out, c0_n7_IO_out, c0_n8_IO_out, c0_n9_IO_out, c0_n10_IO_out, c0_n11_IO_out, c0_n12_IO_out, c0_n13_IO_out, c0_n14_IO_out, c0_n15_IO_out, c0_n16_IO_out, c0_n17_IO_out, c0_n18_IO_out, c0_n19_IO_out, c0_n20_IO_out, c0_n21_IO_out, c0_n22_IO_out, c0_n23_IO_out, c0_n24_IO_out, c0_n25_IO_out, c0_n26_IO_out, c0_n27_IO_out, c0_n28_IO_out, c0_n29_IO_out, c0_n30_IO_out, c0_n31_IO_out, c0_n32_IO_out, c0_n33_IO_out, c0_n34_IO_out, c0_n35_IO_out, c0_n36_IO_out, c0_n37_IO_out, c0_n38_IO_out, c0_n39_IO_out, c0_n40_IO_out, c0_n41_IO_out, c0_n42_IO_out, c0_n43_IO_out, c0_n44_IO_out, c0_n45_IO_out, c0_n46_IO_out, c0_n47_IO_out, c0_n48_IO_out, c0_n49_IO_out, c0_n50_IO_out, c0_n51_IO_out, c0_n52_IO_out, c0_n53_IO_out, c0_n54_IO_out, c0_n55_IO_out, c0_n56_IO_out, c0_n57_IO_out, c0_n58_IO_out, c0_n59_IO_out, c0_n60_IO_out, c0_n61_IO_out, c0_n62_IO_out, c0_n63_IO_out, c0_n64_IO_out, c0_n65_IO_out, c0_n66_IO_out, c0_n67_IO_out, c0_n68_IO_out, c0_n69_IO_out, c0_n70_IO_out, c0_n71_IO_out, c0_n72_IO_out, c0_n73_IO_out, c0_n74_IO_out, c0_n75_IO_out, c0_n76_IO_out, c0_n77_IO_out, c0_n78_IO_out, c0_n79_IO_out, c0_n80_IO_out, c0_n81_IO_out, c0_n82_IO_out, c0_n83_IO_out, c0_n84_IO_out, c0_n85_IO_out, c0_n86_IO_out, c0_n87_IO_out, c0_n88_IO_out, c0_n89_IO_out, c0_n90_IO_out, c0_n91_IO_out, c0_n92_IO_out, c0_n93_IO_out, c0_n94_IO_out, c0_n95_IO_out, c0_n96_IO_out, c0_n97_IO_out, c0_n98_IO_out, c0_n99_IO_out, c0_n100_IO_out, c0_n101_IO_out, c0_n102_IO_out, c0_n103_IO_out, c0_n104_IO_out, c0_n105_IO_out, c0_n106_IO_out, c0_n107_IO_out, c0_n108_IO_out, c0_n109_IO_out, c0_n110_IO_out, c0_n111_IO_out, c0_n112_IO_out, c0_n113_IO_out, c0_n114_IO_out, c0_n115_IO_out, c0_n116_IO_out, c0_n117_IO_out, c0_n118_IO_out, c0_n119_IO_out, c0_n120_IO_out, c0_n121_IO_out, c0_n122_IO_out, c0_n123_IO_out, c0_n124_IO_out, c0_n125_IO_out, c0_n126_IO_out, c0_n127_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c1_n0_IO_out, c1_n1_IO_out, c1_n2_IO_out, c1_n3_IO_out, c1_n4_IO_out, c1_n5_IO_out, c1_n6_IO_out, c1_n7_IO_out, c1_n8_IO_out, c1_n9_IO_out, c1_n10_IO_out, c1_n11_IO_out, c1_n12_IO_out, c1_n13_IO_out, c1_n14_IO_out, c1_n15_IO_out, c1_n16_IO_out, c1_n17_IO_out, c1_n18_IO_out, c1_n19_IO_out, c1_n20_IO_out, c1_n21_IO_out, c1_n22_IO_out, c1_n23_IO_out, c1_n24_IO_out, c1_n25_IO_out, c1_n26_IO_out, c1_n27_IO_out, c1_n28_IO_out, c1_n29_IO_out, c1_n30_IO_out, c1_n31_IO_out, c1_n32_IO_out, c1_n33_IO_out, c1_n34_IO_out, c1_n35_IO_out, c1_n36_IO_out, c1_n37_IO_out, c1_n38_IO_out, c1_n39_IO_out, c1_n40_IO_out, c1_n41_IO_out, c1_n42_IO_out, c1_n43_IO_out, c1_n44_IO_out, c1_n45_IO_out, c1_n46_IO_out, c1_n47_IO_out, c1_n48_IO_out, c1_n49_IO_out, c1_n50_IO_out, c1_n51_IO_out, c1_n52_IO_out, c1_n53_IO_out, c1_n54_IO_out, c1_n55_IO_out, c1_n56_IO_out, c1_n57_IO_out, c1_n58_IO_out, c1_n59_IO_out, c1_n60_IO_out, c1_n61_IO_out, c1_n62_IO_out, c1_n63_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c2_n0_IO_out, c2_n1_IO_out, c2_n2_IO_out, c2_n3_IO_out, c2_n4_IO_out, c2_n5_IO_out, c2_n6_IO_out, c2_n7_IO_out, c2_n8_IO_out, c2_n9_IO_out, c2_n10_IO_out, c2_n11_IO_out, c2_n12_IO_out, c2_n13_IO_out, c2_n14_IO_out, c2_n15_IO_out, c2_n16_IO_out, c2_n17_IO_out, c2_n18_IO_out, c2_n19_IO_out, c2_n20_IO_out, c2_n21_IO_out, c2_n22_IO_out, c2_n23_IO_out, c2_n24_IO_out, c2_n25_IO_out, c2_n26_IO_out, c2_n27_IO_out, c2_n28_IO_out, c2_n29_IO_out, c2_n30_IO_out, c2_n31_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c3_n0_IO_out, c3_n1_IO_out, c3_n2_IO_out, c3_n3_IO_out, c3_n4_IO_out, c3_n5_IO_out, c3_n6_IO_out, c3_n7_IO_out, c3_n8_IO_out, c3_n9_IO_out, c3_n10_IO_out, c3_n11_IO_out, c3_n12_IO_out, c3_n13_IO_out, c3_n14_IO_out, c3_n15_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c4_n0_IO_out, c4_n1_IO_out, c4_n2_IO_out, c4_n3_IO_out, c4_n4_IO_out, c4_n5_IO_out, c4_n6_IO_out, c4_n7_IO_out, c4_n8_IO_out, c4_n9_IO_out, c4_n10_IO_out, c4_n11_IO_out, c4_n12_IO_out, c4_n13_IO_out, c4_n14_IO_out, c4_n15_IO_out, c4_n16_IO_out, c4_n17_IO_out, c4_n18_IO_out, c4_n19_IO_out, c4_n20_IO_out, c4_n21_IO_out, c4_n22_IO_out, c4_n23_IO_out, c4_n24_IO_out, c4_n25_IO_out, c4_n26_IO_out, c4_n27_IO_out, c4_n28_IO_out, c4_n29_IO_out, c4_n30_IO_out, c4_n31_IO_out: SIGNED(BITS -1 DOWNTO 0);
  SIGNAL c5_n0_IO_out, c5_n1_IO_out, c5_n2_IO_out, c5_n3_IO_out, c5_n4_IO_out, c5_n5_IO_out, c5_n6_IO_out, c5_n7_IO_out, c5_n8_IO_out, c5_n9_IO_out, c5_n10_IO_out, c5_n11_IO_out, c5_n12_IO_out, c5_n13_IO_out, c5_n14_IO_out, c5_n15_IO_out, c5_n16_IO_out, c5_n17_IO_out, c5_n18_IO_out, c5_n19_IO_out, c5_n20_IO_out, c5_n21_IO_out, c5_n22_IO_out, c5_n23_IO_out, c5_n24_IO_out, c5_n25_IO_out, c5_n26_IO_out, c5_n27_IO_out, c5_n28_IO_out, c5_n29_IO_out, c5_n30_IO_out, c5_n31_IO_out, c5_n32_IO_out, c5_n33_IO_out, c5_n34_IO_out, c5_n35_IO_out, c5_n36_IO_out, c5_n37_IO_out, c5_n38_IO_out, c5_n39_IO_out, c5_n40_IO_out, c5_n41_IO_out, c5_n42_IO_out, c5_n43_IO_out, c5_n44_IO_out, c5_n45_IO_out, c5_n46_IO_out, c5_n47_IO_out, c5_n48_IO_out, c5_n49_IO_out, c5_n50_IO_out, c5_n51_IO_out, c5_n52_IO_out, c5_n53_IO_out, c5_n54_IO_out, c5_n55_IO_out, c5_n56_IO_out, c5_n57_IO_out, c5_n58_IO_out, c5_n59_IO_out, c5_n60_IO_out, c5_n61_IO_out, c5_n62_IO_out, c5_n63_IO_out: SIGNED(BITS -1 DOWNTO 0);
    SIGNAL reg_IO_in: signed(TOTAL_BITS - 1 DOWNTO 0);
    SIGNAL en_registers: STD_LOGIC;
BEGIN
  en_registers <= update_weights AND clk;
  c1_IO_in <= c0_n0_IO_out & c0_n1_IO_out & c0_n2_IO_out & c0_n3_IO_out & c0_n4_IO_out & c0_n5_IO_out & c0_n6_IO_out & c0_n7_IO_out & c0_n8_IO_out & c0_n9_IO_out & c0_n10_IO_out & c0_n11_IO_out & c0_n12_IO_out & c0_n13_IO_out & c0_n14_IO_out & c0_n15_IO_out & c0_n16_IO_out & c0_n17_IO_out & c0_n18_IO_out & c0_n19_IO_out & c0_n20_IO_out & c0_n21_IO_out & c0_n22_IO_out & c0_n23_IO_out & c0_n24_IO_out & c0_n25_IO_out & c0_n26_IO_out & c0_n27_IO_out & c0_n28_IO_out & c0_n29_IO_out & c0_n30_IO_out & c0_n31_IO_out & c0_n32_IO_out & c0_n33_IO_out & c0_n34_IO_out & c0_n35_IO_out & c0_n36_IO_out & c0_n37_IO_out & c0_n38_IO_out & c0_n39_IO_out & c0_n40_IO_out & c0_n41_IO_out & c0_n42_IO_out & c0_n43_IO_out & c0_n44_IO_out & c0_n45_IO_out & c0_n46_IO_out & c0_n47_IO_out & c0_n48_IO_out & c0_n49_IO_out & c0_n50_IO_out & c0_n51_IO_out & c0_n52_IO_out & c0_n53_IO_out & c0_n54_IO_out & c0_n55_IO_out & c0_n56_IO_out & c0_n57_IO_out & c0_n58_IO_out & c0_n59_IO_out & c0_n60_IO_out & c0_n61_IO_out & c0_n62_IO_out & c0_n63_IO_out & c0_n64_IO_out & c0_n65_IO_out & c0_n66_IO_out & c0_n67_IO_out & c0_n68_IO_out & c0_n69_IO_out & c0_n70_IO_out & c0_n71_IO_out & c0_n72_IO_out & c0_n73_IO_out & c0_n74_IO_out & c0_n75_IO_out & c0_n76_IO_out & c0_n77_IO_out & c0_n78_IO_out & c0_n79_IO_out & c0_n80_IO_out & c0_n81_IO_out & c0_n82_IO_out & c0_n83_IO_out & c0_n84_IO_out & c0_n85_IO_out & c0_n86_IO_out & c0_n87_IO_out & c0_n88_IO_out & c0_n89_IO_out & c0_n90_IO_out & c0_n91_IO_out & c0_n92_IO_out & c0_n93_IO_out & c0_n94_IO_out & c0_n95_IO_out & c0_n96_IO_out & c0_n97_IO_out & c0_n98_IO_out & c0_n99_IO_out & c0_n100_IO_out & c0_n101_IO_out & c0_n102_IO_out & c0_n103_IO_out & c0_n104_IO_out & c0_n105_IO_out & c0_n106_IO_out & c0_n107_IO_out & c0_n108_IO_out & c0_n109_IO_out & c0_n110_IO_out & c0_n111_IO_out & c0_n112_IO_out & c0_n113_IO_out & c0_n114_IO_out & c0_n115_IO_out & c0_n116_IO_out & c0_n117_IO_out & c0_n118_IO_out & c0_n119_IO_out & c0_n120_IO_out & c0_n121_IO_out & c0_n122_IO_out & c0_n123_IO_out & c0_n124_IO_out & c0_n125_IO_out & c0_n126_IO_out & c0_n127_IO_out;
c2_IO_in <= c1_n0_IO_out & c1_n1_IO_out & c1_n2_IO_out & c1_n3_IO_out & c1_n4_IO_out & c1_n5_IO_out & c1_n6_IO_out & c1_n7_IO_out & c1_n8_IO_out & c1_n9_IO_out & c1_n10_IO_out & c1_n11_IO_out & c1_n12_IO_out & c1_n13_IO_out & c1_n14_IO_out & c1_n15_IO_out & c1_n16_IO_out & c1_n17_IO_out & c1_n18_IO_out & c1_n19_IO_out & c1_n20_IO_out & c1_n21_IO_out & c1_n22_IO_out & c1_n23_IO_out & c1_n24_IO_out & c1_n25_IO_out & c1_n26_IO_out & c1_n27_IO_out & c1_n28_IO_out & c1_n29_IO_out & c1_n30_IO_out & c1_n31_IO_out & c1_n32_IO_out & c1_n33_IO_out & c1_n34_IO_out & c1_n35_IO_out & c1_n36_IO_out & c1_n37_IO_out & c1_n38_IO_out & c1_n39_IO_out & c1_n40_IO_out & c1_n41_IO_out & c1_n42_IO_out & c1_n43_IO_out & c1_n44_IO_out & c1_n45_IO_out & c1_n46_IO_out & c1_n47_IO_out & c1_n48_IO_out & c1_n49_IO_out & c1_n50_IO_out & c1_n51_IO_out & c1_n52_IO_out & c1_n53_IO_out & c1_n54_IO_out & c1_n55_IO_out & c1_n56_IO_out & c1_n57_IO_out & c1_n58_IO_out & c1_n59_IO_out & c1_n60_IO_out & c1_n61_IO_out & c1_n62_IO_out & c1_n63_IO_out;
c3_IO_in <= c2_n0_IO_out & c2_n1_IO_out & c2_n2_IO_out & c2_n3_IO_out & c2_n4_IO_out & c2_n5_IO_out & c2_n6_IO_out & c2_n7_IO_out & c2_n8_IO_out & c2_n9_IO_out & c2_n10_IO_out & c2_n11_IO_out & c2_n12_IO_out & c2_n13_IO_out & c2_n14_IO_out & c2_n15_IO_out & c2_n16_IO_out & c2_n17_IO_out & c2_n18_IO_out & c2_n19_IO_out & c2_n20_IO_out & c2_n21_IO_out & c2_n22_IO_out & c2_n23_IO_out & c2_n24_IO_out & c2_n25_IO_out & c2_n26_IO_out & c2_n27_IO_out & c2_n28_IO_out & c2_n29_IO_out & c2_n30_IO_out & c2_n31_IO_out;
c4_IO_in <= c3_n0_IO_out & c3_n1_IO_out & c3_n2_IO_out & c3_n3_IO_out & c3_n4_IO_out & c3_n5_IO_out & c3_n6_IO_out & c3_n7_IO_out & c3_n8_IO_out & c3_n9_IO_out & c3_n10_IO_out & c3_n11_IO_out & c3_n12_IO_out & c3_n13_IO_out & c3_n14_IO_out & c3_n15_IO_out;
c5_IO_in <= c4_n0_IO_out & c4_n1_IO_out & c4_n2_IO_out & c4_n3_IO_out & c4_n4_IO_out & c4_n5_IO_out & c4_n6_IO_out & c4_n7_IO_out & c4_n8_IO_out & c4_n9_IO_out & c4_n10_IO_out & c4_n11_IO_out & c4_n12_IO_out & c4_n13_IO_out & c4_n14_IO_out & c4_n15_IO_out & c4_n16_IO_out & c4_n17_IO_out & c4_n18_IO_out & c4_n19_IO_out & c4_n20_IO_out & c4_n21_IO_out & c4_n22_IO_out & c4_n23_IO_out & c4_n24_IO_out & c4_n25_IO_out & c4_n26_IO_out & c4_n27_IO_out & c4_n28_IO_out & c4_n29_IO_out & c4_n30_IO_out & c4_n31_IO_out;
c6_IO_in <= c5_n0_IO_out & c5_n1_IO_out & c5_n2_IO_out & c5_n3_IO_out & c5_n4_IO_out & c5_n5_IO_out & c5_n6_IO_out & c5_n7_IO_out & c5_n8_IO_out & c5_n9_IO_out & c5_n10_IO_out & c5_n11_IO_out & c5_n12_IO_out & c5_n13_IO_out & c5_n14_IO_out & c5_n15_IO_out & c5_n16_IO_out & c5_n17_IO_out & c5_n18_IO_out & c5_n19_IO_out & c5_n20_IO_out & c5_n21_IO_out & c5_n22_IO_out & c5_n23_IO_out & c5_n24_IO_out & c5_n25_IO_out & c5_n26_IO_out & c5_n27_IO_out & c5_n28_IO_out & c5_n29_IO_out & c5_n30_IO_out & c5_n31_IO_out & c5_n32_IO_out & c5_n33_IO_out & c5_n34_IO_out & c5_n35_IO_out & c5_n36_IO_out & c5_n37_IO_out & c5_n38_IO_out & c5_n39_IO_out & c5_n40_IO_out & c5_n41_IO_out & c5_n42_IO_out & c5_n43_IO_out & c5_n44_IO_out & c5_n45_IO_out & c5_n46_IO_out & c5_n47_IO_out & c5_n48_IO_out & c5_n49_IO_out & c5_n50_IO_out & c5_n51_IO_out & c5_n52_IO_out & c5_n53_IO_out & c5_n54_IO_out & c5_n55_IO_out & c5_n56_IO_out & c5_n57_IO_out & c5_n58_IO_out & c5_n59_IO_out & c5_n60_IO_out & c5_n61_IO_out & c5_n62_IO_out & c5_n63_IO_out;

  PROCESS (clk, rst)
  BEGIN
    IF rst = '1' THEN
      reg_IO_in <= (OTHERS => '0');
    ELSIF clk'event AND clk = '1' THEN
      reg_IO_in <= IO_in;
    END IF;
  END PROCESS;

camada0_inst_0: ENTITY work.camada0_ReLU_128neuron_8bits_784n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> reg_IO_in, 
            c0_n0_W_in=> c0_n0_W_in, 
            c0_n1_W_in=> c0_n1_W_in, 
            c0_n2_W_in=> c0_n2_W_in, 
            c0_n3_W_in=> c0_n3_W_in, 
            c0_n4_W_in=> c0_n4_W_in, 
            c0_n5_W_in=> c0_n5_W_in, 
            c0_n6_W_in=> c0_n6_W_in, 
            c0_n7_W_in=> c0_n7_W_in, 
            c0_n8_W_in=> c0_n8_W_in, 
            c0_n9_W_in=> c0_n9_W_in, 
            c0_n10_W_in=> c0_n10_W_in, 
            c0_n11_W_in=> c0_n11_W_in, 
            c0_n12_W_in=> c0_n12_W_in, 
            c0_n13_W_in=> c0_n13_W_in, 
            c0_n14_W_in=> c0_n14_W_in, 
            c0_n15_W_in=> c0_n15_W_in, 
            c0_n16_W_in=> c0_n16_W_in, 
            c0_n17_W_in=> c0_n17_W_in, 
            c0_n18_W_in=> c0_n18_W_in, 
            c0_n19_W_in=> c0_n19_W_in, 
            c0_n20_W_in=> c0_n20_W_in, 
            c0_n21_W_in=> c0_n21_W_in, 
            c0_n22_W_in=> c0_n22_W_in, 
            c0_n23_W_in=> c0_n23_W_in, 
            c0_n24_W_in=> c0_n24_W_in, 
            c0_n25_W_in=> c0_n25_W_in, 
            c0_n26_W_in=> c0_n26_W_in, 
            c0_n27_W_in=> c0_n27_W_in, 
            c0_n28_W_in=> c0_n28_W_in, 
            c0_n29_W_in=> c0_n29_W_in, 
            c0_n30_W_in=> c0_n30_W_in, 
            c0_n31_W_in=> c0_n31_W_in, 
            c0_n32_W_in=> c0_n32_W_in, 
            c0_n33_W_in=> c0_n33_W_in, 
            c0_n34_W_in=> c0_n34_W_in, 
            c0_n35_W_in=> c0_n35_W_in, 
            c0_n36_W_in=> c0_n36_W_in, 
            c0_n37_W_in=> c0_n37_W_in, 
            c0_n38_W_in=> c0_n38_W_in, 
            c0_n39_W_in=> c0_n39_W_in, 
            c0_n40_W_in=> c0_n40_W_in, 
            c0_n41_W_in=> c0_n41_W_in, 
            c0_n42_W_in=> c0_n42_W_in, 
            c0_n43_W_in=> c0_n43_W_in, 
            c0_n44_W_in=> c0_n44_W_in, 
            c0_n45_W_in=> c0_n45_W_in, 
            c0_n46_W_in=> c0_n46_W_in, 
            c0_n47_W_in=> c0_n47_W_in, 
            c0_n48_W_in=> c0_n48_W_in, 
            c0_n49_W_in=> c0_n49_W_in, 
            c0_n50_W_in=> c0_n50_W_in, 
            c0_n51_W_in=> c0_n51_W_in, 
            c0_n52_W_in=> c0_n52_W_in, 
            c0_n53_W_in=> c0_n53_W_in, 
            c0_n54_W_in=> c0_n54_W_in, 
            c0_n55_W_in=> c0_n55_W_in, 
            c0_n56_W_in=> c0_n56_W_in, 
            c0_n57_W_in=> c0_n57_W_in, 
            c0_n58_W_in=> c0_n58_W_in, 
            c0_n59_W_in=> c0_n59_W_in, 
            c0_n60_W_in=> c0_n60_W_in, 
            c0_n61_W_in=> c0_n61_W_in, 
            c0_n62_W_in=> c0_n62_W_in, 
            c0_n63_W_in=> c0_n63_W_in, 
            c0_n64_W_in=> c0_n64_W_in, 
            c0_n65_W_in=> c0_n65_W_in, 
            c0_n66_W_in=> c0_n66_W_in, 
            c0_n67_W_in=> c0_n67_W_in, 
            c0_n68_W_in=> c0_n68_W_in, 
            c0_n69_W_in=> c0_n69_W_in, 
            c0_n70_W_in=> c0_n70_W_in, 
            c0_n71_W_in=> c0_n71_W_in, 
            c0_n72_W_in=> c0_n72_W_in, 
            c0_n73_W_in=> c0_n73_W_in, 
            c0_n74_W_in=> c0_n74_W_in, 
            c0_n75_W_in=> c0_n75_W_in, 
            c0_n76_W_in=> c0_n76_W_in, 
            c0_n77_W_in=> c0_n77_W_in, 
            c0_n78_W_in=> c0_n78_W_in, 
            c0_n79_W_in=> c0_n79_W_in, 
            c0_n80_W_in=> c0_n80_W_in, 
            c0_n81_W_in=> c0_n81_W_in, 
            c0_n82_W_in=> c0_n82_W_in, 
            c0_n83_W_in=> c0_n83_W_in, 
            c0_n84_W_in=> c0_n84_W_in, 
            c0_n85_W_in=> c0_n85_W_in, 
            c0_n86_W_in=> c0_n86_W_in, 
            c0_n87_W_in=> c0_n87_W_in, 
            c0_n88_W_in=> c0_n88_W_in, 
            c0_n89_W_in=> c0_n89_W_in, 
            c0_n90_W_in=> c0_n90_W_in, 
            c0_n91_W_in=> c0_n91_W_in, 
            c0_n92_W_in=> c0_n92_W_in, 
            c0_n93_W_in=> c0_n93_W_in, 
            c0_n94_W_in=> c0_n94_W_in, 
            c0_n95_W_in=> c0_n95_W_in, 
            c0_n96_W_in=> c0_n96_W_in, 
            c0_n97_W_in=> c0_n97_W_in, 
            c0_n98_W_in=> c0_n98_W_in, 
            c0_n99_W_in=> c0_n99_W_in, 
            c0_n100_W_in=> c0_n100_W_in, 
            c0_n101_W_in=> c0_n101_W_in, 
            c0_n102_W_in=> c0_n102_W_in, 
            c0_n103_W_in=> c0_n103_W_in, 
            c0_n104_W_in=> c0_n104_W_in, 
            c0_n105_W_in=> c0_n105_W_in, 
            c0_n106_W_in=> c0_n106_W_in, 
            c0_n107_W_in=> c0_n107_W_in, 
            c0_n108_W_in=> c0_n108_W_in, 
            c0_n109_W_in=> c0_n109_W_in, 
            c0_n110_W_in=> c0_n110_W_in, 
            c0_n111_W_in=> c0_n111_W_in, 
            c0_n112_W_in=> c0_n112_W_in, 
            c0_n113_W_in=> c0_n113_W_in, 
            c0_n114_W_in=> c0_n114_W_in, 
            c0_n115_W_in=> c0_n115_W_in, 
            c0_n116_W_in=> c0_n116_W_in, 
            c0_n117_W_in=> c0_n117_W_in, 
            c0_n118_W_in=> c0_n118_W_in, 
            c0_n119_W_in=> c0_n119_W_in, 
            c0_n120_W_in=> c0_n120_W_in, 
            c0_n121_W_in=> c0_n121_W_in, 
            c0_n122_W_in=> c0_n122_W_in, 
            c0_n123_W_in=> c0_n123_W_in, 
            c0_n124_W_in=> c0_n124_W_in, 
            c0_n125_W_in=> c0_n125_W_in, 
            c0_n126_W_in=> c0_n126_W_in, 
            c0_n127_W_in=> c0_n127_W_in, 
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c0_n0_IO_out=> c0_n0_IO_out, 
            c0_n1_IO_out=> c0_n1_IO_out, 
            c0_n2_IO_out=> c0_n2_IO_out, 
            c0_n3_IO_out=> c0_n3_IO_out, 
            c0_n4_IO_out=> c0_n4_IO_out, 
            c0_n5_IO_out=> c0_n5_IO_out, 
            c0_n6_IO_out=> c0_n6_IO_out, 
            c0_n7_IO_out=> c0_n7_IO_out, 
            c0_n8_IO_out=> c0_n8_IO_out, 
            c0_n9_IO_out=> c0_n9_IO_out, 
            c0_n10_IO_out=> c0_n10_IO_out, 
            c0_n11_IO_out=> c0_n11_IO_out, 
            c0_n12_IO_out=> c0_n12_IO_out, 
            c0_n13_IO_out=> c0_n13_IO_out, 
            c0_n14_IO_out=> c0_n14_IO_out, 
            c0_n15_IO_out=> c0_n15_IO_out, 
            c0_n16_IO_out=> c0_n16_IO_out, 
            c0_n17_IO_out=> c0_n17_IO_out, 
            c0_n18_IO_out=> c0_n18_IO_out, 
            c0_n19_IO_out=> c0_n19_IO_out, 
            c0_n20_IO_out=> c0_n20_IO_out, 
            c0_n21_IO_out=> c0_n21_IO_out, 
            c0_n22_IO_out=> c0_n22_IO_out, 
            c0_n23_IO_out=> c0_n23_IO_out, 
            c0_n24_IO_out=> c0_n24_IO_out, 
            c0_n25_IO_out=> c0_n25_IO_out, 
            c0_n26_IO_out=> c0_n26_IO_out, 
            c0_n27_IO_out=> c0_n27_IO_out, 
            c0_n28_IO_out=> c0_n28_IO_out, 
            c0_n29_IO_out=> c0_n29_IO_out, 
            c0_n30_IO_out=> c0_n30_IO_out, 
            c0_n31_IO_out=> c0_n31_IO_out, 
            c0_n32_IO_out=> c0_n32_IO_out, 
            c0_n33_IO_out=> c0_n33_IO_out, 
            c0_n34_IO_out=> c0_n34_IO_out, 
            c0_n35_IO_out=> c0_n35_IO_out, 
            c0_n36_IO_out=> c0_n36_IO_out, 
            c0_n37_IO_out=> c0_n37_IO_out, 
            c0_n38_IO_out=> c0_n38_IO_out, 
            c0_n39_IO_out=> c0_n39_IO_out, 
            c0_n40_IO_out=> c0_n40_IO_out, 
            c0_n41_IO_out=> c0_n41_IO_out, 
            c0_n42_IO_out=> c0_n42_IO_out, 
            c0_n43_IO_out=> c0_n43_IO_out, 
            c0_n44_IO_out=> c0_n44_IO_out, 
            c0_n45_IO_out=> c0_n45_IO_out, 
            c0_n46_IO_out=> c0_n46_IO_out, 
            c0_n47_IO_out=> c0_n47_IO_out, 
            c0_n48_IO_out=> c0_n48_IO_out, 
            c0_n49_IO_out=> c0_n49_IO_out, 
            c0_n50_IO_out=> c0_n50_IO_out, 
            c0_n51_IO_out=> c0_n51_IO_out, 
            c0_n52_IO_out=> c0_n52_IO_out, 
            c0_n53_IO_out=> c0_n53_IO_out, 
            c0_n54_IO_out=> c0_n54_IO_out, 
            c0_n55_IO_out=> c0_n55_IO_out, 
            c0_n56_IO_out=> c0_n56_IO_out, 
            c0_n57_IO_out=> c0_n57_IO_out, 
            c0_n58_IO_out=> c0_n58_IO_out, 
            c0_n59_IO_out=> c0_n59_IO_out, 
            c0_n60_IO_out=> c0_n60_IO_out, 
            c0_n61_IO_out=> c0_n61_IO_out, 
            c0_n62_IO_out=> c0_n62_IO_out, 
            c0_n63_IO_out=> c0_n63_IO_out, 
            c0_n64_IO_out=> c0_n64_IO_out, 
            c0_n65_IO_out=> c0_n65_IO_out, 
            c0_n66_IO_out=> c0_n66_IO_out, 
            c0_n67_IO_out=> c0_n67_IO_out, 
            c0_n68_IO_out=> c0_n68_IO_out, 
            c0_n69_IO_out=> c0_n69_IO_out, 
            c0_n70_IO_out=> c0_n70_IO_out, 
            c0_n71_IO_out=> c0_n71_IO_out, 
            c0_n72_IO_out=> c0_n72_IO_out, 
            c0_n73_IO_out=> c0_n73_IO_out, 
            c0_n74_IO_out=> c0_n74_IO_out, 
            c0_n75_IO_out=> c0_n75_IO_out, 
            c0_n76_IO_out=> c0_n76_IO_out, 
            c0_n77_IO_out=> c0_n77_IO_out, 
            c0_n78_IO_out=> c0_n78_IO_out, 
            c0_n79_IO_out=> c0_n79_IO_out, 
            c0_n80_IO_out=> c0_n80_IO_out, 
            c0_n81_IO_out=> c0_n81_IO_out, 
            c0_n82_IO_out=> c0_n82_IO_out, 
            c0_n83_IO_out=> c0_n83_IO_out, 
            c0_n84_IO_out=> c0_n84_IO_out, 
            c0_n85_IO_out=> c0_n85_IO_out, 
            c0_n86_IO_out=> c0_n86_IO_out, 
            c0_n87_IO_out=> c0_n87_IO_out, 
            c0_n88_IO_out=> c0_n88_IO_out, 
            c0_n89_IO_out=> c0_n89_IO_out, 
            c0_n90_IO_out=> c0_n90_IO_out, 
            c0_n91_IO_out=> c0_n91_IO_out, 
            c0_n92_IO_out=> c0_n92_IO_out, 
            c0_n93_IO_out=> c0_n93_IO_out, 
            c0_n94_IO_out=> c0_n94_IO_out, 
            c0_n95_IO_out=> c0_n95_IO_out, 
            c0_n96_IO_out=> c0_n96_IO_out, 
            c0_n97_IO_out=> c0_n97_IO_out, 
            c0_n98_IO_out=> c0_n98_IO_out, 
            c0_n99_IO_out=> c0_n99_IO_out, 
            c0_n100_IO_out=> c0_n100_IO_out, 
            c0_n101_IO_out=> c0_n101_IO_out, 
            c0_n102_IO_out=> c0_n102_IO_out, 
            c0_n103_IO_out=> c0_n103_IO_out, 
            c0_n104_IO_out=> c0_n104_IO_out, 
            c0_n105_IO_out=> c0_n105_IO_out, 
            c0_n106_IO_out=> c0_n106_IO_out, 
            c0_n107_IO_out=> c0_n107_IO_out, 
            c0_n108_IO_out=> c0_n108_IO_out, 
            c0_n109_IO_out=> c0_n109_IO_out, 
            c0_n110_IO_out=> c0_n110_IO_out, 
            c0_n111_IO_out=> c0_n111_IO_out, 
            c0_n112_IO_out=> c0_n112_IO_out, 
            c0_n113_IO_out=> c0_n113_IO_out, 
            c0_n114_IO_out=> c0_n114_IO_out, 
            c0_n115_IO_out=> c0_n115_IO_out, 
            c0_n116_IO_out=> c0_n116_IO_out, 
            c0_n117_IO_out=> c0_n117_IO_out, 
            c0_n118_IO_out=> c0_n118_IO_out, 
            c0_n119_IO_out=> c0_n119_IO_out, 
            c0_n120_IO_out=> c0_n120_IO_out, 
            c0_n121_IO_out=> c0_n121_IO_out, 
            c0_n122_IO_out=> c0_n122_IO_out, 
            c0_n123_IO_out=> c0_n123_IO_out, 
            c0_n124_IO_out=> c0_n124_IO_out, 
            c0_n125_IO_out=> c0_n125_IO_out, 
            c0_n126_IO_out=> c0_n126_IO_out, 
            c0_n127_IO_out=> c0_n127_IO_out, 
            -- ['OUT']['manual'] 
            c0_n0_W_out=> c0_n0_W_out, 
            c0_n1_W_out=> c0_n1_W_out, 
            c0_n2_W_out=> c0_n2_W_out, 
            c0_n3_W_out=> c0_n3_W_out, 
            c0_n4_W_out=> c0_n4_W_out, 
            c0_n5_W_out=> c0_n5_W_out, 
            c0_n6_W_out=> c0_n6_W_out, 
            c0_n7_W_out=> c0_n7_W_out, 
            c0_n8_W_out=> c0_n8_W_out, 
            c0_n9_W_out=> c0_n9_W_out, 
            c0_n10_W_out=> c0_n10_W_out, 
            c0_n11_W_out=> c0_n11_W_out, 
            c0_n12_W_out=> c0_n12_W_out, 
            c0_n13_W_out=> c0_n13_W_out, 
            c0_n14_W_out=> c0_n14_W_out, 
            c0_n15_W_out=> c0_n15_W_out, 
            c0_n16_W_out=> c0_n16_W_out, 
            c0_n17_W_out=> c0_n17_W_out, 
            c0_n18_W_out=> c0_n18_W_out, 
            c0_n19_W_out=> c0_n19_W_out, 
            c0_n20_W_out=> c0_n20_W_out, 
            c0_n21_W_out=> c0_n21_W_out, 
            c0_n22_W_out=> c0_n22_W_out, 
            c0_n23_W_out=> c0_n23_W_out, 
            c0_n24_W_out=> c0_n24_W_out, 
            c0_n25_W_out=> c0_n25_W_out, 
            c0_n26_W_out=> c0_n26_W_out, 
            c0_n27_W_out=> c0_n27_W_out, 
            c0_n28_W_out=> c0_n28_W_out, 
            c0_n29_W_out=> c0_n29_W_out, 
            c0_n30_W_out=> c0_n30_W_out, 
            c0_n31_W_out=> c0_n31_W_out, 
            c0_n32_W_out=> c0_n32_W_out, 
            c0_n33_W_out=> c0_n33_W_out, 
            c0_n34_W_out=> c0_n34_W_out, 
            c0_n35_W_out=> c0_n35_W_out, 
            c0_n36_W_out=> c0_n36_W_out, 
            c0_n37_W_out=> c0_n37_W_out, 
            c0_n38_W_out=> c0_n38_W_out, 
            c0_n39_W_out=> c0_n39_W_out, 
            c0_n40_W_out=> c0_n40_W_out, 
            c0_n41_W_out=> c0_n41_W_out, 
            c0_n42_W_out=> c0_n42_W_out, 
            c0_n43_W_out=> c0_n43_W_out, 
            c0_n44_W_out=> c0_n44_W_out, 
            c0_n45_W_out=> c0_n45_W_out, 
            c0_n46_W_out=> c0_n46_W_out, 
            c0_n47_W_out=> c0_n47_W_out, 
            c0_n48_W_out=> c0_n48_W_out, 
            c0_n49_W_out=> c0_n49_W_out, 
            c0_n50_W_out=> c0_n50_W_out, 
            c0_n51_W_out=> c0_n51_W_out, 
            c0_n52_W_out=> c0_n52_W_out, 
            c0_n53_W_out=> c0_n53_W_out, 
            c0_n54_W_out=> c0_n54_W_out, 
            c0_n55_W_out=> c0_n55_W_out, 
            c0_n56_W_out=> c0_n56_W_out, 
            c0_n57_W_out=> c0_n57_W_out, 
            c0_n58_W_out=> c0_n58_W_out, 
            c0_n59_W_out=> c0_n59_W_out, 
            c0_n60_W_out=> c0_n60_W_out, 
            c0_n61_W_out=> c0_n61_W_out, 
            c0_n62_W_out=> c0_n62_W_out, 
            c0_n63_W_out=> c0_n63_W_out, 
            c0_n64_W_out=> c0_n64_W_out, 
            c0_n65_W_out=> c0_n65_W_out, 
            c0_n66_W_out=> c0_n66_W_out, 
            c0_n67_W_out=> c0_n67_W_out, 
            c0_n68_W_out=> c0_n68_W_out, 
            c0_n69_W_out=> c0_n69_W_out, 
            c0_n70_W_out=> c0_n70_W_out, 
            c0_n71_W_out=> c0_n71_W_out, 
            c0_n72_W_out=> c0_n72_W_out, 
            c0_n73_W_out=> c0_n73_W_out, 
            c0_n74_W_out=> c0_n74_W_out, 
            c0_n75_W_out=> c0_n75_W_out, 
            c0_n76_W_out=> c0_n76_W_out, 
            c0_n77_W_out=> c0_n77_W_out, 
            c0_n78_W_out=> c0_n78_W_out, 
            c0_n79_W_out=> c0_n79_W_out, 
            c0_n80_W_out=> c0_n80_W_out, 
            c0_n81_W_out=> c0_n81_W_out, 
            c0_n82_W_out=> c0_n82_W_out, 
            c0_n83_W_out=> c0_n83_W_out, 
            c0_n84_W_out=> c0_n84_W_out, 
            c0_n85_W_out=> c0_n85_W_out, 
            c0_n86_W_out=> c0_n86_W_out, 
            c0_n87_W_out=> c0_n87_W_out, 
            c0_n88_W_out=> c0_n88_W_out, 
            c0_n89_W_out=> c0_n89_W_out, 
            c0_n90_W_out=> c0_n90_W_out, 
            c0_n91_W_out=> c0_n91_W_out, 
            c0_n92_W_out=> c0_n92_W_out, 
            c0_n93_W_out=> c0_n93_W_out, 
            c0_n94_W_out=> c0_n94_W_out, 
            c0_n95_W_out=> c0_n95_W_out, 
            c0_n96_W_out=> c0_n96_W_out, 
            c0_n97_W_out=> c0_n97_W_out, 
            c0_n98_W_out=> c0_n98_W_out, 
            c0_n99_W_out=> c0_n99_W_out, 
            c0_n100_W_out=> c0_n100_W_out, 
            c0_n101_W_out=> c0_n101_W_out, 
            c0_n102_W_out=> c0_n102_W_out, 
            c0_n103_W_out=> c0_n103_W_out, 
            c0_n104_W_out=> c0_n104_W_out, 
            c0_n105_W_out=> c0_n105_W_out, 
            c0_n106_W_out=> c0_n106_W_out, 
            c0_n107_W_out=> c0_n107_W_out, 
            c0_n108_W_out=> c0_n108_W_out, 
            c0_n109_W_out=> c0_n109_W_out, 
            c0_n110_W_out=> c0_n110_W_out, 
            c0_n111_W_out=> c0_n111_W_out, 
            c0_n112_W_out=> c0_n112_W_out, 
            c0_n113_W_out=> c0_n113_W_out, 
            c0_n114_W_out=> c0_n114_W_out, 
            c0_n115_W_out=> c0_n115_W_out, 
            c0_n116_W_out=> c0_n116_W_out, 
            c0_n117_W_out=> c0_n117_W_out, 
            c0_n118_W_out=> c0_n118_W_out, 
            c0_n119_W_out=> c0_n119_W_out, 
            c0_n120_W_out=> c0_n120_W_out, 
            c0_n121_W_out=> c0_n121_W_out, 
            c0_n122_W_out=> c0_n122_W_out, 
            c0_n123_W_out=> c0_n123_W_out, 
            c0_n124_W_out=> c0_n124_W_out, 
            c0_n125_W_out=> c0_n125_W_out, 
            c0_n126_W_out=> c0_n126_W_out, 
            c0_n127_W_out=> c0_n127_W_out
   );
            
camada1_inst_1: ENTITY work.camada1_ReLU_64neuron_8bits_128n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c1_IO_in, 
            c1_n0_W_in=> c0_n0_W_out,
            c1_n1_W_in=> c0_n1_W_out,
            c1_n2_W_in=> c0_n2_W_out,
            c1_n3_W_in=> c0_n3_W_out,
            c1_n4_W_in=> c0_n4_W_out,
            c1_n5_W_in=> c0_n5_W_out,
            c1_n6_W_in=> c0_n6_W_out,
            c1_n7_W_in=> c0_n7_W_out,
            c1_n8_W_in=> c0_n8_W_out,
            c1_n9_W_in=> c0_n9_W_out,
            c1_n10_W_in=> c0_n10_W_out,
            c1_n11_W_in=> c0_n11_W_out,
            c1_n12_W_in=> c0_n12_W_out,
            c1_n13_W_in=> c0_n13_W_out,
            c1_n14_W_in=> c0_n14_W_out,
            c1_n15_W_in=> c0_n15_W_out,
            c1_n16_W_in=> c0_n16_W_out,
            c1_n17_W_in=> c0_n17_W_out,
            c1_n18_W_in=> c0_n18_W_out,
            c1_n19_W_in=> c0_n19_W_out,
            c1_n20_W_in=> c0_n20_W_out,
            c1_n21_W_in=> c0_n21_W_out,
            c1_n22_W_in=> c0_n22_W_out,
            c1_n23_W_in=> c0_n23_W_out,
            c1_n24_W_in=> c0_n24_W_out,
            c1_n25_W_in=> c0_n25_W_out,
            c1_n26_W_in=> c0_n26_W_out,
            c1_n27_W_in=> c0_n27_W_out,
            c1_n28_W_in=> c0_n28_W_out,
            c1_n29_W_in=> c0_n29_W_out,
            c1_n30_W_in=> c0_n30_W_out,
            c1_n31_W_in=> c0_n31_W_out,
            c1_n32_W_in=> c0_n32_W_out,
            c1_n33_W_in=> c0_n33_W_out,
            c1_n34_W_in=> c0_n34_W_out,
            c1_n35_W_in=> c0_n35_W_out,
            c1_n36_W_in=> c0_n36_W_out,
            c1_n37_W_in=> c0_n37_W_out,
            c1_n38_W_in=> c0_n38_W_out,
            c1_n39_W_in=> c0_n39_W_out,
            c1_n40_W_in=> c0_n40_W_out,
            c1_n41_W_in=> c0_n41_W_out,
            c1_n42_W_in=> c0_n42_W_out,
            c1_n43_W_in=> c0_n43_W_out,
            c1_n44_W_in=> c0_n44_W_out,
            c1_n45_W_in=> c0_n45_W_out,
            c1_n46_W_in=> c0_n46_W_out,
            c1_n47_W_in=> c0_n47_W_out,
            c1_n48_W_in=> c0_n48_W_out,
            c1_n49_W_in=> c0_n49_W_out,
            c1_n50_W_in=> c0_n50_W_out,
            c1_n51_W_in=> c0_n51_W_out,
            c1_n52_W_in=> c0_n52_W_out,
            c1_n53_W_in=> c0_n53_W_out,
            c1_n54_W_in=> c0_n54_W_out,
            c1_n55_W_in=> c0_n55_W_out,
            c1_n56_W_in=> c0_n56_W_out,
            c1_n57_W_in=> c0_n57_W_out,
            c1_n58_W_in=> c0_n58_W_out,
            c1_n59_W_in=> c0_n59_W_out,
            c1_n60_W_in=> c0_n60_W_out,
            c1_n61_W_in=> c0_n61_W_out,
            c1_n62_W_in=> c0_n62_W_out,
            c1_n63_W_in=> c0_n63_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c1_n0_IO_out=> c1_n0_IO_out, 
            c1_n1_IO_out=> c1_n1_IO_out, 
            c1_n2_IO_out=> c1_n2_IO_out, 
            c1_n3_IO_out=> c1_n3_IO_out, 
            c1_n4_IO_out=> c1_n4_IO_out, 
            c1_n5_IO_out=> c1_n5_IO_out, 
            c1_n6_IO_out=> c1_n6_IO_out, 
            c1_n7_IO_out=> c1_n7_IO_out, 
            c1_n8_IO_out=> c1_n8_IO_out, 
            c1_n9_IO_out=> c1_n9_IO_out, 
            c1_n10_IO_out=> c1_n10_IO_out, 
            c1_n11_IO_out=> c1_n11_IO_out, 
            c1_n12_IO_out=> c1_n12_IO_out, 
            c1_n13_IO_out=> c1_n13_IO_out, 
            c1_n14_IO_out=> c1_n14_IO_out, 
            c1_n15_IO_out=> c1_n15_IO_out, 
            c1_n16_IO_out=> c1_n16_IO_out, 
            c1_n17_IO_out=> c1_n17_IO_out, 
            c1_n18_IO_out=> c1_n18_IO_out, 
            c1_n19_IO_out=> c1_n19_IO_out, 
            c1_n20_IO_out=> c1_n20_IO_out, 
            c1_n21_IO_out=> c1_n21_IO_out, 
            c1_n22_IO_out=> c1_n22_IO_out, 
            c1_n23_IO_out=> c1_n23_IO_out, 
            c1_n24_IO_out=> c1_n24_IO_out, 
            c1_n25_IO_out=> c1_n25_IO_out, 
            c1_n26_IO_out=> c1_n26_IO_out, 
            c1_n27_IO_out=> c1_n27_IO_out, 
            c1_n28_IO_out=> c1_n28_IO_out, 
            c1_n29_IO_out=> c1_n29_IO_out, 
            c1_n30_IO_out=> c1_n30_IO_out, 
            c1_n31_IO_out=> c1_n31_IO_out, 
            c1_n32_IO_out=> c1_n32_IO_out, 
            c1_n33_IO_out=> c1_n33_IO_out, 
            c1_n34_IO_out=> c1_n34_IO_out, 
            c1_n35_IO_out=> c1_n35_IO_out, 
            c1_n36_IO_out=> c1_n36_IO_out, 
            c1_n37_IO_out=> c1_n37_IO_out, 
            c1_n38_IO_out=> c1_n38_IO_out, 
            c1_n39_IO_out=> c1_n39_IO_out, 
            c1_n40_IO_out=> c1_n40_IO_out, 
            c1_n41_IO_out=> c1_n41_IO_out, 
            c1_n42_IO_out=> c1_n42_IO_out, 
            c1_n43_IO_out=> c1_n43_IO_out, 
            c1_n44_IO_out=> c1_n44_IO_out, 
            c1_n45_IO_out=> c1_n45_IO_out, 
            c1_n46_IO_out=> c1_n46_IO_out, 
            c1_n47_IO_out=> c1_n47_IO_out, 
            c1_n48_IO_out=> c1_n48_IO_out, 
            c1_n49_IO_out=> c1_n49_IO_out, 
            c1_n50_IO_out=> c1_n50_IO_out, 
            c1_n51_IO_out=> c1_n51_IO_out, 
            c1_n52_IO_out=> c1_n52_IO_out, 
            c1_n53_IO_out=> c1_n53_IO_out, 
            c1_n54_IO_out=> c1_n54_IO_out, 
            c1_n55_IO_out=> c1_n55_IO_out, 
            c1_n56_IO_out=> c1_n56_IO_out, 
            c1_n57_IO_out=> c1_n57_IO_out, 
            c1_n58_IO_out=> c1_n58_IO_out, 
            c1_n59_IO_out=> c1_n59_IO_out, 
            c1_n60_IO_out=> c1_n60_IO_out, 
            c1_n61_IO_out=> c1_n61_IO_out, 
            c1_n62_IO_out=> c1_n62_IO_out, 
            c1_n63_IO_out=> c1_n63_IO_out, 
            -- ['OUT']['manual'] 
            c1_n0_W_out=> c1_n0_W_out, 
            c1_n1_W_out=> c1_n1_W_out, 
            c1_n2_W_out=> c1_n2_W_out, 
            c1_n3_W_out=> c1_n3_W_out, 
            c1_n4_W_out=> c1_n4_W_out, 
            c1_n5_W_out=> c1_n5_W_out, 
            c1_n6_W_out=> c1_n6_W_out, 
            c1_n7_W_out=> c1_n7_W_out, 
            c1_n8_W_out=> c1_n8_W_out, 
            c1_n9_W_out=> c1_n9_W_out, 
            c1_n10_W_out=> c1_n10_W_out, 
            c1_n11_W_out=> c1_n11_W_out, 
            c1_n12_W_out=> c1_n12_W_out, 
            c1_n13_W_out=> c1_n13_W_out, 
            c1_n14_W_out=> c1_n14_W_out, 
            c1_n15_W_out=> c1_n15_W_out, 
            c1_n16_W_out=> c1_n16_W_out, 
            c1_n17_W_out=> c1_n17_W_out, 
            c1_n18_W_out=> c1_n18_W_out, 
            c1_n19_W_out=> c1_n19_W_out, 
            c1_n20_W_out=> c1_n20_W_out, 
            c1_n21_W_out=> c1_n21_W_out, 
            c1_n22_W_out=> c1_n22_W_out, 
            c1_n23_W_out=> c1_n23_W_out, 
            c1_n24_W_out=> c1_n24_W_out, 
            c1_n25_W_out=> c1_n25_W_out, 
            c1_n26_W_out=> c1_n26_W_out, 
            c1_n27_W_out=> c1_n27_W_out, 
            c1_n28_W_out=> c1_n28_W_out, 
            c1_n29_W_out=> c1_n29_W_out, 
            c1_n30_W_out=> c1_n30_W_out, 
            c1_n31_W_out=> c1_n31_W_out, 
            c1_n32_W_out=> c1_n32_W_out, 
            c1_n33_W_out=> c1_n33_W_out, 
            c1_n34_W_out=> c1_n34_W_out, 
            c1_n35_W_out=> c1_n35_W_out, 
            c1_n36_W_out=> c1_n36_W_out, 
            c1_n37_W_out=> c1_n37_W_out, 
            c1_n38_W_out=> c1_n38_W_out, 
            c1_n39_W_out=> c1_n39_W_out, 
            c1_n40_W_out=> c1_n40_W_out, 
            c1_n41_W_out=> c1_n41_W_out, 
            c1_n42_W_out=> c1_n42_W_out, 
            c1_n43_W_out=> c1_n43_W_out, 
            c1_n44_W_out=> c1_n44_W_out, 
            c1_n45_W_out=> c1_n45_W_out, 
            c1_n46_W_out=> c1_n46_W_out, 
            c1_n47_W_out=> c1_n47_W_out, 
            c1_n48_W_out=> c1_n48_W_out, 
            c1_n49_W_out=> c1_n49_W_out, 
            c1_n50_W_out=> c1_n50_W_out, 
            c1_n51_W_out=> c1_n51_W_out, 
            c1_n52_W_out=> c1_n52_W_out, 
            c1_n53_W_out=> c1_n53_W_out, 
            c1_n54_W_out=> c1_n54_W_out, 
            c1_n55_W_out=> c1_n55_W_out, 
            c1_n56_W_out=> c1_n56_W_out, 
            c1_n57_W_out=> c1_n57_W_out, 
            c1_n58_W_out=> c1_n58_W_out, 
            c1_n59_W_out=> c1_n59_W_out, 
            c1_n60_W_out=> c1_n60_W_out, 
            c1_n61_W_out=> c1_n61_W_out, 
            c1_n62_W_out=> c1_n62_W_out, 
            c1_n63_W_out=> c1_n63_W_out
   );
            
camada2_inst_2: ENTITY work.camada2_ReLU_32neuron_8bits_64n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c2_IO_in, 
            c2_n0_W_in=> c1_n0_W_out,
            c2_n1_W_in=> c1_n1_W_out,
            c2_n2_W_in=> c1_n2_W_out,
            c2_n3_W_in=> c1_n3_W_out,
            c2_n4_W_in=> c1_n4_W_out,
            c2_n5_W_in=> c1_n5_W_out,
            c2_n6_W_in=> c1_n6_W_out,
            c2_n7_W_in=> c1_n7_W_out,
            c2_n8_W_in=> c1_n8_W_out,
            c2_n9_W_in=> c1_n9_W_out,
            c2_n10_W_in=> c1_n10_W_out,
            c2_n11_W_in=> c1_n11_W_out,
            c2_n12_W_in=> c1_n12_W_out,
            c2_n13_W_in=> c1_n13_W_out,
            c2_n14_W_in=> c1_n14_W_out,
            c2_n15_W_in=> c1_n15_W_out,
            c2_n16_W_in=> c1_n16_W_out,
            c2_n17_W_in=> c1_n17_W_out,
            c2_n18_W_in=> c1_n18_W_out,
            c2_n19_W_in=> c1_n19_W_out,
            c2_n20_W_in=> c1_n20_W_out,
            c2_n21_W_in=> c1_n21_W_out,
            c2_n22_W_in=> c1_n22_W_out,
            c2_n23_W_in=> c1_n23_W_out,
            c2_n24_W_in=> c1_n24_W_out,
            c2_n25_W_in=> c1_n25_W_out,
            c2_n26_W_in=> c1_n26_W_out,
            c2_n27_W_in=> c1_n27_W_out,
            c2_n28_W_in=> c1_n28_W_out,
            c2_n29_W_in=> c1_n29_W_out,
            c2_n30_W_in=> c1_n30_W_out,
            c2_n31_W_in=> c1_n31_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c2_n0_IO_out=> c2_n0_IO_out, 
            c2_n1_IO_out=> c2_n1_IO_out, 
            c2_n2_IO_out=> c2_n2_IO_out, 
            c2_n3_IO_out=> c2_n3_IO_out, 
            c2_n4_IO_out=> c2_n4_IO_out, 
            c2_n5_IO_out=> c2_n5_IO_out, 
            c2_n6_IO_out=> c2_n6_IO_out, 
            c2_n7_IO_out=> c2_n7_IO_out, 
            c2_n8_IO_out=> c2_n8_IO_out, 
            c2_n9_IO_out=> c2_n9_IO_out, 
            c2_n10_IO_out=> c2_n10_IO_out, 
            c2_n11_IO_out=> c2_n11_IO_out, 
            c2_n12_IO_out=> c2_n12_IO_out, 
            c2_n13_IO_out=> c2_n13_IO_out, 
            c2_n14_IO_out=> c2_n14_IO_out, 
            c2_n15_IO_out=> c2_n15_IO_out, 
            c2_n16_IO_out=> c2_n16_IO_out, 
            c2_n17_IO_out=> c2_n17_IO_out, 
            c2_n18_IO_out=> c2_n18_IO_out, 
            c2_n19_IO_out=> c2_n19_IO_out, 
            c2_n20_IO_out=> c2_n20_IO_out, 
            c2_n21_IO_out=> c2_n21_IO_out, 
            c2_n22_IO_out=> c2_n22_IO_out, 
            c2_n23_IO_out=> c2_n23_IO_out, 
            c2_n24_IO_out=> c2_n24_IO_out, 
            c2_n25_IO_out=> c2_n25_IO_out, 
            c2_n26_IO_out=> c2_n26_IO_out, 
            c2_n27_IO_out=> c2_n27_IO_out, 
            c2_n28_IO_out=> c2_n28_IO_out, 
            c2_n29_IO_out=> c2_n29_IO_out, 
            c2_n30_IO_out=> c2_n30_IO_out, 
            c2_n31_IO_out=> c2_n31_IO_out, 
            -- ['OUT']['manual'] 
            c2_n0_W_out=> c2_n0_W_out, 
            c2_n1_W_out=> c2_n1_W_out, 
            c2_n2_W_out=> c2_n2_W_out, 
            c2_n3_W_out=> c2_n3_W_out, 
            c2_n4_W_out=> c2_n4_W_out, 
            c2_n5_W_out=> c2_n5_W_out, 
            c2_n6_W_out=> c2_n6_W_out, 
            c2_n7_W_out=> c2_n7_W_out, 
            c2_n8_W_out=> c2_n8_W_out, 
            c2_n9_W_out=> c2_n9_W_out, 
            c2_n10_W_out=> c2_n10_W_out, 
            c2_n11_W_out=> c2_n11_W_out, 
            c2_n12_W_out=> c2_n12_W_out, 
            c2_n13_W_out=> c2_n13_W_out, 
            c2_n14_W_out=> c2_n14_W_out, 
            c2_n15_W_out=> c2_n15_W_out, 
            c2_n16_W_out=> c2_n16_W_out, 
            c2_n17_W_out=> c2_n17_W_out, 
            c2_n18_W_out=> c2_n18_W_out, 
            c2_n19_W_out=> c2_n19_W_out, 
            c2_n20_W_out=> c2_n20_W_out, 
            c2_n21_W_out=> c2_n21_W_out, 
            c2_n22_W_out=> c2_n22_W_out, 
            c2_n23_W_out=> c2_n23_W_out, 
            c2_n24_W_out=> c2_n24_W_out, 
            c2_n25_W_out=> c2_n25_W_out, 
            c2_n26_W_out=> c2_n26_W_out, 
            c2_n27_W_out=> c2_n27_W_out, 
            c2_n28_W_out=> c2_n28_W_out, 
            c2_n29_W_out=> c2_n29_W_out, 
            c2_n30_W_out=> c2_n30_W_out, 
            c2_n31_W_out=> c2_n31_W_out
   );
            
camada3_inst_3: ENTITY work.camada3_ReLU_16neuron_8bits_32n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c3_IO_in, 
            c3_n0_W_in=> c2_n0_W_out,
            c3_n1_W_in=> c2_n1_W_out,
            c3_n2_W_in=> c2_n2_W_out,
            c3_n3_W_in=> c2_n3_W_out,
            c3_n4_W_in=> c2_n4_W_out,
            c3_n5_W_in=> c2_n5_W_out,
            c3_n6_W_in=> c2_n6_W_out,
            c3_n7_W_in=> c2_n7_W_out,
            c3_n8_W_in=> c2_n8_W_out,
            c3_n9_W_in=> c2_n9_W_out,
            c3_n10_W_in=> c2_n10_W_out,
            c3_n11_W_in=> c2_n11_W_out,
            c3_n12_W_in=> c2_n12_W_out,
            c3_n13_W_in=> c2_n13_W_out,
            c3_n14_W_in=> c2_n14_W_out,
            c3_n15_W_in=> c2_n15_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c3_n0_IO_out=> c3_n0_IO_out, 
            c3_n1_IO_out=> c3_n1_IO_out, 
            c3_n2_IO_out=> c3_n2_IO_out, 
            c3_n3_IO_out=> c3_n3_IO_out, 
            c3_n4_IO_out=> c3_n4_IO_out, 
            c3_n5_IO_out=> c3_n5_IO_out, 
            c3_n6_IO_out=> c3_n6_IO_out, 
            c3_n7_IO_out=> c3_n7_IO_out, 
            c3_n8_IO_out=> c3_n8_IO_out, 
            c3_n9_IO_out=> c3_n9_IO_out, 
            c3_n10_IO_out=> c3_n10_IO_out, 
            c3_n11_IO_out=> c3_n11_IO_out, 
            c3_n12_IO_out=> c3_n12_IO_out, 
            c3_n13_IO_out=> c3_n13_IO_out, 
            c3_n14_IO_out=> c3_n14_IO_out, 
            c3_n15_IO_out=> c3_n15_IO_out, 
            -- ['OUT']['manual'] 
            c3_n0_W_out=> c3_n0_W_out, 
            c3_n1_W_out=> c3_n1_W_out, 
            c3_n2_W_out=> c3_n2_W_out, 
            c3_n3_W_out=> c3_n3_W_out, 
            c3_n4_W_out=> c3_n4_W_out, 
            c3_n5_W_out=> c3_n5_W_out, 
            c3_n6_W_out=> c3_n6_W_out, 
            c3_n7_W_out=> c3_n7_W_out, 
            c3_n8_W_out=> c3_n8_W_out, 
            c3_n9_W_out=> c3_n9_W_out, 
            c3_n10_W_out=> c3_n10_W_out, 
            c3_n11_W_out=> c3_n11_W_out, 
            c3_n12_W_out=> c3_n12_W_out, 
            c3_n13_W_out=> c3_n13_W_out, 
            c3_n14_W_out=> c3_n14_W_out, 
            c3_n15_W_out=> c3_n15_W_out
   );
            
camada4_inst_4: ENTITY work.camada4_ReLU_32neuron_8bits_16n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c4_IO_in, 
            c4_n0_W_in=> c3_n0_W_out,
            c4_n1_W_in=> c3_n1_W_out,
            c4_n2_W_in=> c3_n2_W_out,
            c4_n3_W_in=> c3_n3_W_out,
            c4_n4_W_in=> c3_n4_W_out,
            c4_n5_W_in=> c3_n5_W_out,
            c4_n6_W_in=> c3_n6_W_out,
            c4_n7_W_in=> c3_n7_W_out,
            c4_n8_W_in=> c3_n8_W_out,
            c4_n9_W_in=> c3_n9_W_out,
            c4_n10_W_in=> c3_n10_W_out,
            c4_n11_W_in=> c3_n11_W_out,
            c4_n12_W_in=> c3_n12_W_out,
            c4_n13_W_in=> c3_n13_W_out,
            c4_n14_W_in=> c3_n14_W_out,
            c4_n15_W_in=> c3_n15_W_out,
            c4_n16_W_in=> c2_n16_W_out,
            c4_n17_W_in=> c2_n17_W_out,
            c4_n18_W_in=> c2_n18_W_out,
            c4_n19_W_in=> c2_n19_W_out,
            c4_n20_W_in=> c2_n20_W_out,
            c4_n21_W_in=> c2_n21_W_out,
            c4_n22_W_in=> c2_n22_W_out,
            c4_n23_W_in=> c2_n23_W_out,
            c4_n24_W_in=> c2_n24_W_out,
            c4_n25_W_in=> c2_n25_W_out,
            c4_n26_W_in=> c2_n26_W_out,
            c4_n27_W_in=> c2_n27_W_out,
            c4_n28_W_in=> c2_n28_W_out,
            c4_n29_W_in=> c2_n29_W_out,
            c4_n30_W_in=> c2_n30_W_out,
            c4_n31_W_in=> c2_n31_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c4_n0_IO_out=> c4_n0_IO_out, 
            c4_n1_IO_out=> c4_n1_IO_out, 
            c4_n2_IO_out=> c4_n2_IO_out, 
            c4_n3_IO_out=> c4_n3_IO_out, 
            c4_n4_IO_out=> c4_n4_IO_out, 
            c4_n5_IO_out=> c4_n5_IO_out, 
            c4_n6_IO_out=> c4_n6_IO_out, 
            c4_n7_IO_out=> c4_n7_IO_out, 
            c4_n8_IO_out=> c4_n8_IO_out, 
            c4_n9_IO_out=> c4_n9_IO_out, 
            c4_n10_IO_out=> c4_n10_IO_out, 
            c4_n11_IO_out=> c4_n11_IO_out, 
            c4_n12_IO_out=> c4_n12_IO_out, 
            c4_n13_IO_out=> c4_n13_IO_out, 
            c4_n14_IO_out=> c4_n14_IO_out, 
            c4_n15_IO_out=> c4_n15_IO_out, 
            c4_n16_IO_out=> c4_n16_IO_out, 
            c4_n17_IO_out=> c4_n17_IO_out, 
            c4_n18_IO_out=> c4_n18_IO_out, 
            c4_n19_IO_out=> c4_n19_IO_out, 
            c4_n20_IO_out=> c4_n20_IO_out, 
            c4_n21_IO_out=> c4_n21_IO_out, 
            c4_n22_IO_out=> c4_n22_IO_out, 
            c4_n23_IO_out=> c4_n23_IO_out, 
            c4_n24_IO_out=> c4_n24_IO_out, 
            c4_n25_IO_out=> c4_n25_IO_out, 
            c4_n26_IO_out=> c4_n26_IO_out, 
            c4_n27_IO_out=> c4_n27_IO_out, 
            c4_n28_IO_out=> c4_n28_IO_out, 
            c4_n29_IO_out=> c4_n29_IO_out, 
            c4_n30_IO_out=> c4_n30_IO_out, 
            c4_n31_IO_out=> c4_n31_IO_out, 
            -- ['OUT']['manual'] 
            c4_n0_W_out=> c4_n0_W_out, 
            c4_n1_W_out=> c4_n1_W_out, 
            c4_n2_W_out=> c4_n2_W_out, 
            c4_n3_W_out=> c4_n3_W_out, 
            c4_n4_W_out=> c4_n4_W_out, 
            c4_n5_W_out=> c4_n5_W_out, 
            c4_n6_W_out=> c4_n6_W_out, 
            c4_n7_W_out=> c4_n7_W_out, 
            c4_n8_W_out=> c4_n8_W_out, 
            c4_n9_W_out=> c4_n9_W_out, 
            c4_n10_W_out=> c4_n10_W_out, 
            c4_n11_W_out=> c4_n11_W_out, 
            c4_n12_W_out=> c4_n12_W_out, 
            c4_n13_W_out=> c4_n13_W_out, 
            c4_n14_W_out=> c4_n14_W_out, 
            c4_n15_W_out=> c4_n15_W_out, 
            c4_n16_W_out=> c4_n16_W_out, 
            c4_n17_W_out=> c4_n17_W_out, 
            c4_n18_W_out=> c4_n18_W_out, 
            c4_n19_W_out=> c4_n19_W_out, 
            c4_n20_W_out=> c4_n20_W_out, 
            c4_n21_W_out=> c4_n21_W_out, 
            c4_n22_W_out=> c4_n22_W_out, 
            c4_n23_W_out=> c4_n23_W_out, 
            c4_n24_W_out=> c4_n24_W_out, 
            c4_n25_W_out=> c4_n25_W_out, 
            c4_n26_W_out=> c4_n26_W_out, 
            c4_n27_W_out=> c4_n27_W_out, 
            c4_n28_W_out=> c4_n28_W_out, 
            c4_n29_W_out=> c4_n29_W_out, 
            c4_n30_W_out=> c4_n30_W_out, 
            c4_n31_W_out=> c4_n31_W_out
   );
            
camada5_inst_5: ENTITY work.camada5_ReLU_64neuron_8bits_32n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c5_IO_in, 
            c5_n0_W_in=> c4_n0_W_out,
            c5_n1_W_in=> c4_n1_W_out,
            c5_n2_W_in=> c4_n2_W_out,
            c5_n3_W_in=> c4_n3_W_out,
            c5_n4_W_in=> c4_n4_W_out,
            c5_n5_W_in=> c4_n5_W_out,
            c5_n6_W_in=> c4_n6_W_out,
            c5_n7_W_in=> c4_n7_W_out,
            c5_n8_W_in=> c4_n8_W_out,
            c5_n9_W_in=> c4_n9_W_out,
            c5_n10_W_in=> c4_n10_W_out,
            c5_n11_W_in=> c4_n11_W_out,
            c5_n12_W_in=> c4_n12_W_out,
            c5_n13_W_in=> c4_n13_W_out,
            c5_n14_W_in=> c4_n14_W_out,
            c5_n15_W_in=> c4_n15_W_out,
            c5_n16_W_in=> c4_n16_W_out,
            c5_n17_W_in=> c4_n17_W_out,
            c5_n18_W_in=> c4_n18_W_out,
            c5_n19_W_in=> c4_n19_W_out,
            c5_n20_W_in=> c4_n20_W_out,
            c5_n21_W_in=> c4_n21_W_out,
            c5_n22_W_in=> c4_n22_W_out,
            c5_n23_W_in=> c4_n23_W_out,
            c5_n24_W_in=> c4_n24_W_out,
            c5_n25_W_in=> c4_n25_W_out,
            c5_n26_W_in=> c4_n26_W_out,
            c5_n27_W_in=> c4_n27_W_out,
            c5_n28_W_in=> c4_n28_W_out,
            c5_n29_W_in=> c4_n29_W_out,
            c5_n30_W_in=> c4_n30_W_out,
            c5_n31_W_in=> c4_n31_W_out,
            c5_n32_W_in=> c1_n32_W_out,
            c5_n33_W_in=> c1_n33_W_out,
            c5_n34_W_in=> c1_n34_W_out,
            c5_n35_W_in=> c1_n35_W_out,
            c5_n36_W_in=> c1_n36_W_out,
            c5_n37_W_in=> c1_n37_W_out,
            c5_n38_W_in=> c1_n38_W_out,
            c5_n39_W_in=> c1_n39_W_out,
            c5_n40_W_in=> c1_n40_W_out,
            c5_n41_W_in=> c1_n41_W_out,
            c5_n42_W_in=> c1_n42_W_out,
            c5_n43_W_in=> c1_n43_W_out,
            c5_n44_W_in=> c1_n44_W_out,
            c5_n45_W_in=> c1_n45_W_out,
            c5_n46_W_in=> c1_n46_W_out,
            c5_n47_W_in=> c1_n47_W_out,
            c5_n48_W_in=> c1_n48_W_out,
            c5_n49_W_in=> c1_n49_W_out,
            c5_n50_W_in=> c1_n50_W_out,
            c5_n51_W_in=> c1_n51_W_out,
            c5_n52_W_in=> c1_n52_W_out,
            c5_n53_W_in=> c1_n53_W_out,
            c5_n54_W_in=> c1_n54_W_out,
            c5_n55_W_in=> c1_n55_W_out,
            c5_n56_W_in=> c1_n56_W_out,
            c5_n57_W_in=> c1_n57_W_out,
            c5_n58_W_in=> c1_n58_W_out,
            c5_n59_W_in=> c1_n59_W_out,
            c5_n60_W_in=> c1_n60_W_out,
            c5_n61_W_in=> c1_n61_W_out,
            c5_n62_W_in=> c1_n62_W_out,
            c5_n63_W_in=> c1_n63_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c5_n0_IO_out=> c5_n0_IO_out, 
            c5_n1_IO_out=> c5_n1_IO_out, 
            c5_n2_IO_out=> c5_n2_IO_out, 
            c5_n3_IO_out=> c5_n3_IO_out, 
            c5_n4_IO_out=> c5_n4_IO_out, 
            c5_n5_IO_out=> c5_n5_IO_out, 
            c5_n6_IO_out=> c5_n6_IO_out, 
            c5_n7_IO_out=> c5_n7_IO_out, 
            c5_n8_IO_out=> c5_n8_IO_out, 
            c5_n9_IO_out=> c5_n9_IO_out, 
            c5_n10_IO_out=> c5_n10_IO_out, 
            c5_n11_IO_out=> c5_n11_IO_out, 
            c5_n12_IO_out=> c5_n12_IO_out, 
            c5_n13_IO_out=> c5_n13_IO_out, 
            c5_n14_IO_out=> c5_n14_IO_out, 
            c5_n15_IO_out=> c5_n15_IO_out, 
            c5_n16_IO_out=> c5_n16_IO_out, 
            c5_n17_IO_out=> c5_n17_IO_out, 
            c5_n18_IO_out=> c5_n18_IO_out, 
            c5_n19_IO_out=> c5_n19_IO_out, 
            c5_n20_IO_out=> c5_n20_IO_out, 
            c5_n21_IO_out=> c5_n21_IO_out, 
            c5_n22_IO_out=> c5_n22_IO_out, 
            c5_n23_IO_out=> c5_n23_IO_out, 
            c5_n24_IO_out=> c5_n24_IO_out, 
            c5_n25_IO_out=> c5_n25_IO_out, 
            c5_n26_IO_out=> c5_n26_IO_out, 
            c5_n27_IO_out=> c5_n27_IO_out, 
            c5_n28_IO_out=> c5_n28_IO_out, 
            c5_n29_IO_out=> c5_n29_IO_out, 
            c5_n30_IO_out=> c5_n30_IO_out, 
            c5_n31_IO_out=> c5_n31_IO_out, 
            c5_n32_IO_out=> c5_n32_IO_out, 
            c5_n33_IO_out=> c5_n33_IO_out, 
            c5_n34_IO_out=> c5_n34_IO_out, 
            c5_n35_IO_out=> c5_n35_IO_out, 
            c5_n36_IO_out=> c5_n36_IO_out, 
            c5_n37_IO_out=> c5_n37_IO_out, 
            c5_n38_IO_out=> c5_n38_IO_out, 
            c5_n39_IO_out=> c5_n39_IO_out, 
            c5_n40_IO_out=> c5_n40_IO_out, 
            c5_n41_IO_out=> c5_n41_IO_out, 
            c5_n42_IO_out=> c5_n42_IO_out, 
            c5_n43_IO_out=> c5_n43_IO_out, 
            c5_n44_IO_out=> c5_n44_IO_out, 
            c5_n45_IO_out=> c5_n45_IO_out, 
            c5_n46_IO_out=> c5_n46_IO_out, 
            c5_n47_IO_out=> c5_n47_IO_out, 
            c5_n48_IO_out=> c5_n48_IO_out, 
            c5_n49_IO_out=> c5_n49_IO_out, 
            c5_n50_IO_out=> c5_n50_IO_out, 
            c5_n51_IO_out=> c5_n51_IO_out, 
            c5_n52_IO_out=> c5_n52_IO_out, 
            c5_n53_IO_out=> c5_n53_IO_out, 
            c5_n54_IO_out=> c5_n54_IO_out, 
            c5_n55_IO_out=> c5_n55_IO_out, 
            c5_n56_IO_out=> c5_n56_IO_out, 
            c5_n57_IO_out=> c5_n57_IO_out, 
            c5_n58_IO_out=> c5_n58_IO_out, 
            c5_n59_IO_out=> c5_n59_IO_out, 
            c5_n60_IO_out=> c5_n60_IO_out, 
            c5_n61_IO_out=> c5_n61_IO_out, 
            c5_n62_IO_out=> c5_n62_IO_out, 
            c5_n63_IO_out=> c5_n63_IO_out, 
            -- ['OUT']['manual'] 
            c5_n0_W_out=> c5_n0_W_out, 
            c5_n1_W_out=> c5_n1_W_out, 
            c5_n2_W_out=> c5_n2_W_out, 
            c5_n3_W_out=> c5_n3_W_out, 
            c5_n4_W_out=> c5_n4_W_out, 
            c5_n5_W_out=> c5_n5_W_out, 
            c5_n6_W_out=> c5_n6_W_out, 
            c5_n7_W_out=> c5_n7_W_out, 
            c5_n8_W_out=> c5_n8_W_out, 
            c5_n9_W_out=> c5_n9_W_out, 
            c5_n10_W_out=> c5_n10_W_out, 
            c5_n11_W_out=> c5_n11_W_out, 
            c5_n12_W_out=> c5_n12_W_out, 
            c5_n13_W_out=> c5_n13_W_out, 
            c5_n14_W_out=> c5_n14_W_out, 
            c5_n15_W_out=> c5_n15_W_out, 
            c5_n16_W_out=> c5_n16_W_out, 
            c5_n17_W_out=> c5_n17_W_out, 
            c5_n18_W_out=> c5_n18_W_out, 
            c5_n19_W_out=> c5_n19_W_out, 
            c5_n20_W_out=> c5_n20_W_out, 
            c5_n21_W_out=> c5_n21_W_out, 
            c5_n22_W_out=> c5_n22_W_out, 
            c5_n23_W_out=> c5_n23_W_out, 
            c5_n24_W_out=> c5_n24_W_out, 
            c5_n25_W_out=> c5_n25_W_out, 
            c5_n26_W_out=> c5_n26_W_out, 
            c5_n27_W_out=> c5_n27_W_out, 
            c5_n28_W_out=> c5_n28_W_out, 
            c5_n29_W_out=> c5_n29_W_out, 
            c5_n30_W_out=> c5_n30_W_out, 
            c5_n31_W_out=> c5_n31_W_out, 
            c5_n32_W_out=> c5_n32_W_out, 
            c5_n33_W_out=> c5_n33_W_out, 
            c5_n34_W_out=> c5_n34_W_out, 
            c5_n35_W_out=> c5_n35_W_out, 
            c5_n36_W_out=> c5_n36_W_out, 
            c5_n37_W_out=> c5_n37_W_out, 
            c5_n38_W_out=> c5_n38_W_out, 
            c5_n39_W_out=> c5_n39_W_out, 
            c5_n40_W_out=> c5_n40_W_out, 
            c5_n41_W_out=> c5_n41_W_out, 
            c5_n42_W_out=> c5_n42_W_out, 
            c5_n43_W_out=> c5_n43_W_out, 
            c5_n44_W_out=> c5_n44_W_out, 
            c5_n45_W_out=> c5_n45_W_out, 
            c5_n46_W_out=> c5_n46_W_out, 
            c5_n47_W_out=> c5_n47_W_out, 
            c5_n48_W_out=> c5_n48_W_out, 
            c5_n49_W_out=> c5_n49_W_out, 
            c5_n50_W_out=> c5_n50_W_out, 
            c5_n51_W_out=> c5_n51_W_out, 
            c5_n52_W_out=> c5_n52_W_out, 
            c5_n53_W_out=> c5_n53_W_out, 
            c5_n54_W_out=> c5_n54_W_out, 
            c5_n55_W_out=> c5_n55_W_out, 
            c5_n56_W_out=> c5_n56_W_out, 
            c5_n57_W_out=> c5_n57_W_out, 
            c5_n58_W_out=> c5_n58_W_out, 
            c5_n59_W_out=> c5_n59_W_out, 
            c5_n60_W_out=> c5_n60_W_out, 
            c5_n61_W_out=> c5_n61_W_out, 
            c5_n62_W_out=> c5_n62_W_out, 
            c5_n63_W_out=> c5_n63_W_out
   );
            
camada6_inst_6: ENTITY work.camada6_Sigmoid_128neuron_8bits_64n_signed
   PORT MAP (
            ---------- Entradas ----------
            -- ['IN']['STD_LOGIC'] 
            clk=> clk, 
            rst=> rst, 
            update_weights=> en_registers, 
            -- ['IN']['manual'] 
            IO_in=> c6_IO_in, 
            c6_n0_W_in=> c5_n0_W_out,
            c6_n1_W_in=> c5_n1_W_out,
            c6_n2_W_in=> c5_n2_W_out,
            c6_n3_W_in=> c5_n3_W_out,
            c6_n4_W_in=> c5_n4_W_out,
            c6_n5_W_in=> c5_n5_W_out,
            c6_n6_W_in=> c5_n6_W_out,
            c6_n7_W_in=> c5_n7_W_out,
            c6_n8_W_in=> c5_n8_W_out,
            c6_n9_W_in=> c5_n9_W_out,
            c6_n10_W_in=> c5_n10_W_out,
            c6_n11_W_in=> c5_n11_W_out,
            c6_n12_W_in=> c5_n12_W_out,
            c6_n13_W_in=> c5_n13_W_out,
            c6_n14_W_in=> c5_n14_W_out,
            c6_n15_W_in=> c5_n15_W_out,
            c6_n16_W_in=> c5_n16_W_out,
            c6_n17_W_in=> c5_n17_W_out,
            c6_n18_W_in=> c5_n18_W_out,
            c6_n19_W_in=> c5_n19_W_out,
            c6_n20_W_in=> c5_n20_W_out,
            c6_n21_W_in=> c5_n21_W_out,
            c6_n22_W_in=> c5_n22_W_out,
            c6_n23_W_in=> c5_n23_W_out,
            c6_n24_W_in=> c5_n24_W_out,
            c6_n25_W_in=> c5_n25_W_out,
            c6_n26_W_in=> c5_n26_W_out,
            c6_n27_W_in=> c5_n27_W_out,
            c6_n28_W_in=> c5_n28_W_out,
            c6_n29_W_in=> c5_n29_W_out,
            c6_n30_W_in=> c5_n30_W_out,
            c6_n31_W_in=> c5_n31_W_out,
            c6_n32_W_in=> c5_n32_W_out,
            c6_n33_W_in=> c5_n33_W_out,
            c6_n34_W_in=> c5_n34_W_out,
            c6_n35_W_in=> c5_n35_W_out,
            c6_n36_W_in=> c5_n36_W_out,
            c6_n37_W_in=> c5_n37_W_out,
            c6_n38_W_in=> c5_n38_W_out,
            c6_n39_W_in=> c5_n39_W_out,
            c6_n40_W_in=> c5_n40_W_out,
            c6_n41_W_in=> c5_n41_W_out,
            c6_n42_W_in=> c5_n42_W_out,
            c6_n43_W_in=> c5_n43_W_out,
            c6_n44_W_in=> c5_n44_W_out,
            c6_n45_W_in=> c5_n45_W_out,
            c6_n46_W_in=> c5_n46_W_out,
            c6_n47_W_in=> c5_n47_W_out,
            c6_n48_W_in=> c5_n48_W_out,
            c6_n49_W_in=> c5_n49_W_out,
            c6_n50_W_in=> c5_n50_W_out,
            c6_n51_W_in=> c5_n51_W_out,
            c6_n52_W_in=> c5_n52_W_out,
            c6_n53_W_in=> c5_n53_W_out,
            c6_n54_W_in=> c5_n54_W_out,
            c6_n55_W_in=> c5_n55_W_out,
            c6_n56_W_in=> c5_n56_W_out,
            c6_n57_W_in=> c5_n57_W_out,
            c6_n58_W_in=> c5_n58_W_out,
            c6_n59_W_in=> c5_n59_W_out,
            c6_n60_W_in=> c5_n60_W_out,
            c6_n61_W_in=> c5_n61_W_out,
            c6_n62_W_in=> c5_n62_W_out,
            c6_n63_W_in=> c5_n63_W_out,
            c6_n64_W_in=> c0_n64_W_out,
            c6_n65_W_in=> c0_n65_W_out,
            c6_n66_W_in=> c0_n66_W_out,
            c6_n67_W_in=> c0_n67_W_out,
            c6_n68_W_in=> c0_n68_W_out,
            c6_n69_W_in=> c0_n69_W_out,
            c6_n70_W_in=> c0_n70_W_out,
            c6_n71_W_in=> c0_n71_W_out,
            c6_n72_W_in=> c0_n72_W_out,
            c6_n73_W_in=> c0_n73_W_out,
            c6_n74_W_in=> c0_n74_W_out,
            c6_n75_W_in=> c0_n75_W_out,
            c6_n76_W_in=> c0_n76_W_out,
            c6_n77_W_in=> c0_n77_W_out,
            c6_n78_W_in=> c0_n78_W_out,
            c6_n79_W_in=> c0_n79_W_out,
            c6_n80_W_in=> c0_n80_W_out,
            c6_n81_W_in=> c0_n81_W_out,
            c6_n82_W_in=> c0_n82_W_out,
            c6_n83_W_in=> c0_n83_W_out,
            c6_n84_W_in=> c0_n84_W_out,
            c6_n85_W_in=> c0_n85_W_out,
            c6_n86_W_in=> c0_n86_W_out,
            c6_n87_W_in=> c0_n87_W_out,
            c6_n88_W_in=> c0_n88_W_out,
            c6_n89_W_in=> c0_n89_W_out,
            c6_n90_W_in=> c0_n90_W_out,
            c6_n91_W_in=> c0_n91_W_out,
            c6_n92_W_in=> c0_n92_W_out,
            c6_n93_W_in=> c0_n93_W_out,
            c6_n94_W_in=> c0_n94_W_out,
            c6_n95_W_in=> c0_n95_W_out,
            c6_n96_W_in=> c0_n96_W_out,
            c6_n97_W_in=> c0_n97_W_out,
            c6_n98_W_in=> c0_n98_W_out,
            c6_n99_W_in=> c0_n99_W_out,
            c6_n100_W_in=> c0_n100_W_out,
            c6_n101_W_in=> c0_n101_W_out,
            c6_n102_W_in=> c0_n102_W_out,
            c6_n103_W_in=> c0_n103_W_out,
            c6_n104_W_in=> c0_n104_W_out,
            c6_n105_W_in=> c0_n105_W_out,
            c6_n106_W_in=> c0_n106_W_out,
            c6_n107_W_in=> c0_n107_W_out,
            c6_n108_W_in=> c0_n108_W_out,
            c6_n109_W_in=> c0_n109_W_out,
            c6_n110_W_in=> c0_n110_W_out,
            c6_n111_W_in=> c0_n111_W_out,
            c6_n112_W_in=> c0_n112_W_out,
            c6_n113_W_in=> c0_n113_W_out,
            c6_n114_W_in=> c0_n114_W_out,
            c6_n115_W_in=> c0_n115_W_out,
            c6_n116_W_in=> c0_n116_W_out,
            c6_n117_W_in=> c0_n117_W_out,
            c6_n118_W_in=> c0_n118_W_out,
            c6_n119_W_in=> c0_n119_W_out,
            c6_n120_W_in=> c0_n120_W_out,
            c6_n121_W_in=> c0_n121_W_out,
            c6_n122_W_in=> c0_n122_W_out,
            c6_n123_W_in=> c0_n123_W_out,
            c6_n124_W_in=> c0_n124_W_out,
            c6_n125_W_in=> c0_n125_W_out,
            c6_n126_W_in=> c0_n126_W_out,
            c6_n127_W_in=> c0_n127_W_out,
            ---------- Saidas ----------
            -- ['OUT']['SIGNED'] 
            c6_n0_IO_out=> c6_n0_IO_out, 
            c6_n1_IO_out=> c6_n1_IO_out, 
            c6_n2_IO_out=> c6_n2_IO_out, 
            c6_n3_IO_out=> c6_n3_IO_out, 
            c6_n4_IO_out=> c6_n4_IO_out, 
            c6_n5_IO_out=> c6_n5_IO_out, 
            c6_n6_IO_out=> c6_n6_IO_out, 
            c6_n7_IO_out=> c6_n7_IO_out, 
            c6_n8_IO_out=> c6_n8_IO_out, 
            c6_n9_IO_out=> c6_n9_IO_out, 
            c6_n10_IO_out=> c6_n10_IO_out, 
            c6_n11_IO_out=> c6_n11_IO_out, 
            c6_n12_IO_out=> c6_n12_IO_out, 
            c6_n13_IO_out=> c6_n13_IO_out, 
            c6_n14_IO_out=> c6_n14_IO_out, 
            c6_n15_IO_out=> c6_n15_IO_out, 
            c6_n16_IO_out=> c6_n16_IO_out, 
            c6_n17_IO_out=> c6_n17_IO_out, 
            c6_n18_IO_out=> c6_n18_IO_out, 
            c6_n19_IO_out=> c6_n19_IO_out, 
            c6_n20_IO_out=> c6_n20_IO_out, 
            c6_n21_IO_out=> c6_n21_IO_out, 
            c6_n22_IO_out=> c6_n22_IO_out, 
            c6_n23_IO_out=> c6_n23_IO_out, 
            c6_n24_IO_out=> c6_n24_IO_out, 
            c6_n25_IO_out=> c6_n25_IO_out, 
            c6_n26_IO_out=> c6_n26_IO_out, 
            c6_n27_IO_out=> c6_n27_IO_out, 
            c6_n28_IO_out=> c6_n28_IO_out, 
            c6_n29_IO_out=> c6_n29_IO_out, 
            c6_n30_IO_out=> c6_n30_IO_out, 
            c6_n31_IO_out=> c6_n31_IO_out, 
            c6_n32_IO_out=> c6_n32_IO_out, 
            c6_n33_IO_out=> c6_n33_IO_out, 
            c6_n34_IO_out=> c6_n34_IO_out, 
            c6_n35_IO_out=> c6_n35_IO_out, 
            c6_n36_IO_out=> c6_n36_IO_out, 
            c6_n37_IO_out=> c6_n37_IO_out, 
            c6_n38_IO_out=> c6_n38_IO_out, 
            c6_n39_IO_out=> c6_n39_IO_out, 
            c6_n40_IO_out=> c6_n40_IO_out, 
            c6_n41_IO_out=> c6_n41_IO_out, 
            c6_n42_IO_out=> c6_n42_IO_out, 
            c6_n43_IO_out=> c6_n43_IO_out, 
            c6_n44_IO_out=> c6_n44_IO_out, 
            c6_n45_IO_out=> c6_n45_IO_out, 
            c6_n46_IO_out=> c6_n46_IO_out, 
            c6_n47_IO_out=> c6_n47_IO_out, 
            c6_n48_IO_out=> c6_n48_IO_out, 
            c6_n49_IO_out=> c6_n49_IO_out, 
            c6_n50_IO_out=> c6_n50_IO_out, 
            c6_n51_IO_out=> c6_n51_IO_out, 
            c6_n52_IO_out=> c6_n52_IO_out, 
            c6_n53_IO_out=> c6_n53_IO_out, 
            c6_n54_IO_out=> c6_n54_IO_out, 
            c6_n55_IO_out=> c6_n55_IO_out, 
            c6_n56_IO_out=> c6_n56_IO_out, 
            c6_n57_IO_out=> c6_n57_IO_out, 
            c6_n58_IO_out=> c6_n58_IO_out, 
            c6_n59_IO_out=> c6_n59_IO_out, 
            c6_n60_IO_out=> c6_n60_IO_out, 
            c6_n61_IO_out=> c6_n61_IO_out, 
            c6_n62_IO_out=> c6_n62_IO_out, 
            c6_n63_IO_out=> c6_n63_IO_out, 
            c6_n64_IO_out=> c6_n64_IO_out, 
            c6_n65_IO_out=> c6_n65_IO_out, 
            c6_n66_IO_out=> c6_n66_IO_out, 
            c6_n67_IO_out=> c6_n67_IO_out, 
            c6_n68_IO_out=> c6_n68_IO_out, 
            c6_n69_IO_out=> c6_n69_IO_out, 
            c6_n70_IO_out=> c6_n70_IO_out, 
            c6_n71_IO_out=> c6_n71_IO_out, 
            c6_n72_IO_out=> c6_n72_IO_out, 
            c6_n73_IO_out=> c6_n73_IO_out, 
            c6_n74_IO_out=> c6_n74_IO_out, 
            c6_n75_IO_out=> c6_n75_IO_out, 
            c6_n76_IO_out=> c6_n76_IO_out, 
            c6_n77_IO_out=> c6_n77_IO_out, 
            c6_n78_IO_out=> c6_n78_IO_out, 
            c6_n79_IO_out=> c6_n79_IO_out, 
            c6_n80_IO_out=> c6_n80_IO_out, 
            c6_n81_IO_out=> c6_n81_IO_out, 
            c6_n82_IO_out=> c6_n82_IO_out, 
            c6_n83_IO_out=> c6_n83_IO_out, 
            c6_n84_IO_out=> c6_n84_IO_out, 
            c6_n85_IO_out=> c6_n85_IO_out, 
            c6_n86_IO_out=> c6_n86_IO_out, 
            c6_n87_IO_out=> c6_n87_IO_out, 
            c6_n88_IO_out=> c6_n88_IO_out, 
            c6_n89_IO_out=> c6_n89_IO_out, 
            c6_n90_IO_out=> c6_n90_IO_out, 
            c6_n91_IO_out=> c6_n91_IO_out, 
            c6_n92_IO_out=> c6_n92_IO_out, 
            c6_n93_IO_out=> c6_n93_IO_out, 
            c6_n94_IO_out=> c6_n94_IO_out, 
            c6_n95_IO_out=> c6_n95_IO_out, 
            c6_n96_IO_out=> c6_n96_IO_out, 
            c6_n97_IO_out=> c6_n97_IO_out, 
            c6_n98_IO_out=> c6_n98_IO_out, 
            c6_n99_IO_out=> c6_n99_IO_out, 
            c6_n100_IO_out=> c6_n100_IO_out, 
            c6_n101_IO_out=> c6_n101_IO_out, 
            c6_n102_IO_out=> c6_n102_IO_out, 
            c6_n103_IO_out=> c6_n103_IO_out, 
            c6_n104_IO_out=> c6_n104_IO_out, 
            c6_n105_IO_out=> c6_n105_IO_out, 
            c6_n106_IO_out=> c6_n106_IO_out, 
            c6_n107_IO_out=> c6_n107_IO_out, 
            c6_n108_IO_out=> c6_n108_IO_out, 
            c6_n109_IO_out=> c6_n109_IO_out, 
            c6_n110_IO_out=> c6_n110_IO_out, 
            c6_n111_IO_out=> c6_n111_IO_out, 
            c6_n112_IO_out=> c6_n112_IO_out, 
            c6_n113_IO_out=> c6_n113_IO_out, 
            c6_n114_IO_out=> c6_n114_IO_out, 
            c6_n115_IO_out=> c6_n115_IO_out, 
            c6_n116_IO_out=> c6_n116_IO_out, 
            c6_n117_IO_out=> c6_n117_IO_out, 
            c6_n118_IO_out=> c6_n118_IO_out, 
            c6_n119_IO_out=> c6_n119_IO_out, 
            c6_n120_IO_out=> c6_n120_IO_out, 
            c6_n121_IO_out=> c6_n121_IO_out, 
            c6_n122_IO_out=> c6_n122_IO_out, 
            c6_n123_IO_out=> c6_n123_IO_out, 
            c6_n124_IO_out=> c6_n124_IO_out, 
            c6_n125_IO_out=> c6_n125_IO_out, 
            c6_n126_IO_out=> c6_n126_IO_out, 
            c6_n127_IO_out=> c6_n127_IO_out
   );
            
END ARCHITECTURE;
